----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07.11.2022 19:01:24
-- Design Name: 
-- Module Name: layer_template - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity layer is
    Port ( 
        x : in STD_LOGIC_VECTOR;
        y : out STD_LOGIC_VECTOR
   );
end layer;

architecture layer_1 of layer is

    Component perceptron
    Generic (
        WEIGHTS : STD_LOGIC_VECTOR;
        SHIFT : Integer;     -- number of shift (left + or right -)
        B : Integer;          -- bias of batch norm
        BATCH_POSITIVE : Boolean    
    );
    Port ( 
        x : in STD_LOGIC_VECTOR;
        y : out STD_LOGIC_VECTOR
   );
    end component;
    
    -- Signals
    signal p0_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p0_out : STD_LOGIC;
	signal p1_in : STD_LOGIC_VECTOR(0 to 59 - 1);
	signal p1_out : STD_LOGIC;
	signal p2_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p2_out : STD_LOGIC;
	signal p3_in : STD_LOGIC_VECTOR(0 to 13 - 1);
	signal p3_out : STD_LOGIC;
	signal p4_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p4_out : STD_LOGIC;
	signal p5_in : STD_LOGIC_VECTOR(0 to 59 - 1);
	signal p5_out : STD_LOGIC;
	signal p6_in : STD_LOGIC_VECTOR(0 to 44 - 1);
	signal p6_out : STD_LOGIC;
	signal p7_in : STD_LOGIC_VECTOR(0 to 53 - 1);
	signal p7_out : STD_LOGIC;
	signal p8_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p8_out : STD_LOGIC;
	signal p9_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p9_out : STD_LOGIC;
	signal p10_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p10_out : STD_LOGIC;
	signal p11_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p11_out : STD_LOGIC;
	signal p12_in : STD_LOGIC_VECTOR(0 to 62 - 1);
	signal p12_out : STD_LOGIC;
	signal p13_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p13_out : STD_LOGIC;
	signal p14_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p14_out : STD_LOGIC;
	signal p15_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p15_out : STD_LOGIC;
	signal p16_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p16_out : STD_LOGIC;
	signal p17_in : STD_LOGIC_VECTOR(0 to 65 - 1);
	signal p17_out : STD_LOGIC;
	signal p18_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p18_out : STD_LOGIC;
	signal p19_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p19_out : STD_LOGIC;
	signal p20_in : STD_LOGIC_VECTOR(0 to 70 - 1);
	signal p20_out : STD_LOGIC;
	signal p21_in : STD_LOGIC_VECTOR(0 to 55 - 1);
	signal p21_out : STD_LOGIC;
	signal p22_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p22_out : STD_LOGIC;
	signal p23_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p23_out : STD_LOGIC;
	signal p24_in : STD_LOGIC_VECTOR(0 to 65 - 1);
	signal p24_out : STD_LOGIC;
	signal p25_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p25_out : STD_LOGIC;
	signal p26_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p26_out : STD_LOGIC;
	signal p27_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p27_out : STD_LOGIC;
	signal p28_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p28_out : STD_LOGIC;
	signal p29_in : STD_LOGIC_VECTOR(0 to 63 - 1);
	signal p29_out : STD_LOGIC;
	signal p30_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p30_out : STD_LOGIC;
	signal p31_in : STD_LOGIC_VECTOR(0 to 85 - 1);
	signal p31_out : STD_LOGIC;
	signal p32_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p32_out : STD_LOGIC;
	signal p33_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p33_out : STD_LOGIC;
	signal p34_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p34_out : STD_LOGIC;
	signal p35_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p35_out : STD_LOGIC;
	signal p36_in : STD_LOGIC_VECTOR(0 to 67 - 1);
	signal p36_out : STD_LOGIC;
	signal p37_in : STD_LOGIC_VECTOR(0 to 48 - 1);
	signal p37_out : STD_LOGIC;
	signal p38_in : STD_LOGIC_VECTOR(0 to 45 - 1);
	signal p38_out : STD_LOGIC;
	signal p39_in : STD_LOGIC_VECTOR(0 to 56 - 1);
	signal p39_out : STD_LOGIC;
	signal p40_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p40_out : STD_LOGIC;
	signal p41_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p41_out : STD_LOGIC;
	signal p42_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p42_out : STD_LOGIC;
	signal p43_in : STD_LOGIC_VECTOR(0 to 86 - 1);
	signal p43_out : STD_LOGIC;
	signal p44_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p44_out : STD_LOGIC;
	signal p45_in : STD_LOGIC_VECTOR(0 to 64 - 1);
	signal p45_out : STD_LOGIC;
	signal p46_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p46_out : STD_LOGIC;
	signal p47_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p47_out : STD_LOGIC;
	signal p48_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p48_out : STD_LOGIC;
	signal p49_in : STD_LOGIC_VECTOR(0 to 69 - 1);
	signal p49_out : STD_LOGIC;
	signal p50_in : STD_LOGIC_VECTOR(0 to 47 - 1);
	signal p50_out : STD_LOGIC;
	signal p51_in : STD_LOGIC_VECTOR(0 to 51 - 1);
	signal p51_out : STD_LOGIC;
	signal p52_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p52_out : STD_LOGIC;
	signal p53_in : STD_LOGIC_VECTOR(0 to 45 - 1);
	signal p53_out : STD_LOGIC;
	signal p54_in : STD_LOGIC_VECTOR(0 to 47 - 1);
	signal p54_out : STD_LOGIC;
	signal p55_in : STD_LOGIC_VECTOR(0 to 57 - 1);
	signal p55_out : STD_LOGIC;
	signal p56_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p56_out : STD_LOGIC;
	signal p57_in : STD_LOGIC_VECTOR(0 to 64 - 1);
	signal p57_out : STD_LOGIC;
	signal p58_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p58_out : STD_LOGIC;
	signal p59_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p59_out : STD_LOGIC;
	signal p60_in : STD_LOGIC_VECTOR(0 to 52 - 1);
	signal p60_out : STD_LOGIC;
	signal p61_in : STD_LOGIC_VECTOR(0 to 71 - 1);
	signal p61_out : STD_LOGIC;
	signal p62_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p62_out : STD_LOGIC;
	signal p63_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p63_out : STD_LOGIC;
	signal p64_in : STD_LOGIC_VECTOR(0 to 54 - 1);
	signal p64_out : STD_LOGIC;
	signal p65_in : STD_LOGIC_VECTOR(0 to 44 - 1);
	signal p65_out : STD_LOGIC;
	signal p66_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p66_out : STD_LOGIC;
	signal p67_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p67_out : STD_LOGIC;
	signal p68_in : STD_LOGIC_VECTOR(0 to 54 - 1);
	signal p68_out : STD_LOGIC;
	signal p69_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p69_out : STD_LOGIC;
	signal p70_in : STD_LOGIC_VECTOR(0 to 59 - 1);
	signal p70_out : STD_LOGIC;
	signal p71_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p71_out : STD_LOGIC;
	signal p72_in : STD_LOGIC_VECTOR(0 to 45 - 1);
	signal p72_out : STD_LOGIC;
	signal p73_in : STD_LOGIC_VECTOR(0 to 53 - 1);
	signal p73_out : STD_LOGIC;
	signal p74_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p74_out : STD_LOGIC;
	signal p75_in : STD_LOGIC_VECTOR(0 to 59 - 1);
	signal p75_out : STD_LOGIC;
	signal p76_in : STD_LOGIC_VECTOR(0 to 56 - 1);
	signal p76_out : STD_LOGIC;
	signal p77_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p77_out : STD_LOGIC;
	signal p78_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p78_out : STD_LOGIC;
	signal p79_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p79_out : STD_LOGIC;
	signal p80_in : STD_LOGIC_VECTOR(0 to 57 - 1);
	signal p80_out : STD_LOGIC;
	signal p81_in : STD_LOGIC_VECTOR(0 to 45 - 1);
	signal p81_out : STD_LOGIC;
	signal p82_in : STD_LOGIC_VECTOR(0 to 55 - 1);
	signal p82_out : STD_LOGIC;
	signal p83_in : STD_LOGIC_VECTOR(0 to 48 - 1);
	signal p83_out : STD_LOGIC;
	signal p84_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p84_out : STD_LOGIC;
	signal p85_in : STD_LOGIC_VECTOR(0 to 52 - 1);
	signal p85_out : STD_LOGIC;
	signal p86_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p86_out : STD_LOGIC;
	signal p87_in : STD_LOGIC_VECTOR(0 to 50 - 1);
	signal p87_out : STD_LOGIC;
	signal p88_in : STD_LOGIC_VECTOR(0 to 50 - 1);
	signal p88_out : STD_LOGIC;
	signal p89_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p89_out : STD_LOGIC;
	signal p90_in : STD_LOGIC_VECTOR(0 to 58 - 1);
	signal p90_out : STD_LOGIC;
	signal p91_in : STD_LOGIC_VECTOR(0 to 60 - 1);
	signal p91_out : STD_LOGIC;
	signal p92_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p92_out : STD_LOGIC;
	signal p93_in : STD_LOGIC_VECTOR(0 to 45 - 1);
	signal p93_out : STD_LOGIC;
	signal p94_in : STD_LOGIC_VECTOR(0 to 44 - 1);
	signal p94_out : STD_LOGIC;
	signal p95_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p95_out : STD_LOGIC;
	signal p96_in : STD_LOGIC_VECTOR(0 to 80 - 1);
	signal p96_out : STD_LOGIC;
	signal p97_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p97_out : STD_LOGIC;
	signal p98_in : STD_LOGIC_VECTOR(0 to 64 - 1);
	signal p98_out : STD_LOGIC;
	signal p99_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p99_out : STD_LOGIC;
	signal p100_in : STD_LOGIC_VECTOR(0 to 51 - 1);
	signal p100_out : STD_LOGIC;
	signal p101_in : STD_LOGIC_VECTOR(0 to 71 - 1);
	signal p101_out : STD_LOGIC;
	signal p102_in : STD_LOGIC_VECTOR(0 to 49 - 1);
	signal p102_out : STD_LOGIC;
	signal p103_in : STD_LOGIC_VECTOR(0 to 14 - 1);
	signal p103_out : STD_LOGIC;
	signal p104_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p104_out : STD_LOGIC;
	signal p105_in : STD_LOGIC_VECTOR(0 to 51 - 1);
	signal p105_out : STD_LOGIC;
	signal p106_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p106_out : STD_LOGIC;
	signal p107_in : STD_LOGIC_VECTOR(0 to 49 - 1);
	signal p107_out : STD_LOGIC;
	signal p108_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p108_out : STD_LOGIC;
	signal p109_in : STD_LOGIC_VECTOR(0 to 72 - 1);
	signal p109_out : STD_LOGIC;
	signal p110_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p110_out : STD_LOGIC;
	signal p111_in : STD_LOGIC_VECTOR(0 to 57 - 1);
	signal p111_out : STD_LOGIC;
	signal p112_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p112_out : STD_LOGIC;
	signal p113_in : STD_LOGIC_VECTOR(0 to 57 - 1);
	signal p113_out : STD_LOGIC;
	signal p114_in : STD_LOGIC_VECTOR(0 to 49 - 1);
	signal p114_out : STD_LOGIC;
	signal p115_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p115_out : STD_LOGIC;
	signal p116_in : STD_LOGIC_VECTOR(0 to 74 - 1);
	signal p116_out : STD_LOGIC;
	signal p117_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p117_out : STD_LOGIC;
	signal p118_in : STD_LOGIC_VECTOR(0 to 44 - 1);
	signal p118_out : STD_LOGIC;
	signal p119_in : STD_LOGIC_VECTOR(0 to 50 - 1);
	signal p119_out : STD_LOGIC;
	signal p120_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p120_out : STD_LOGIC;
	signal p121_in : STD_LOGIC_VECTOR(0 to 65 - 1);
	signal p121_out : STD_LOGIC;
	signal p122_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p122_out : STD_LOGIC;
	signal p123_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p123_out : STD_LOGIC;
	signal p124_in : STD_LOGIC_VECTOR(0 to 46 - 1);
	signal p124_out : STD_LOGIC;
	signal p125_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p125_out : STD_LOGIC;
	signal p126_in : STD_LOGIC_VECTOR(0 to 65 - 1);
	signal p126_out : STD_LOGIC;
	signal p127_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p127_out : STD_LOGIC;
	signal p128_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p128_out : STD_LOGIC;
	signal p129_in : STD_LOGIC_VECTOR(0 to 46 - 1);
	signal p129_out : STD_LOGIC;
	signal p130_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p130_out : STD_LOGIC;
	signal p131_in : STD_LOGIC_VECTOR(0 to 54 - 1);
	signal p131_out : STD_LOGIC;
	signal p132_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p132_out : STD_LOGIC;
	signal p133_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p133_out : STD_LOGIC;
	signal p134_in : STD_LOGIC_VECTOR(0 to 53 - 1);
	signal p134_out : STD_LOGIC;
	signal p135_in : STD_LOGIC_VECTOR(0 to 71 - 1);
	signal p135_out : STD_LOGIC;
	signal p136_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p136_out : STD_LOGIC;
	signal p137_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p137_out : STD_LOGIC;
	signal p138_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p138_out : STD_LOGIC;
	signal p139_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p139_out : STD_LOGIC;
	signal p140_in : STD_LOGIC_VECTOR(0 to 55 - 1);
	signal p140_out : STD_LOGIC;
	signal p141_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p141_out : STD_LOGIC;
	signal p142_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p142_out : STD_LOGIC;
	signal p143_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p143_out : STD_LOGIC;
	signal p144_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p144_out : STD_LOGIC;
	signal p145_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p145_out : STD_LOGIC;
	signal p146_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p146_out : STD_LOGIC;
	signal p147_in : STD_LOGIC_VECTOR(0 to 69 - 1);
	signal p147_out : STD_LOGIC;
	signal p148_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p148_out : STD_LOGIC;
	signal p149_in : STD_LOGIC_VECTOR(0 to 54 - 1);
	signal p149_out : STD_LOGIC;
	signal p150_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p150_out : STD_LOGIC;
	signal p151_in : STD_LOGIC_VECTOR(0 to 46 - 1);
	signal p151_out : STD_LOGIC;
	signal p152_in : STD_LOGIC_VECTOR(0 to 71 - 1);
	signal p152_out : STD_LOGIC;
	signal p153_in : STD_LOGIC_VECTOR(0 to 68 - 1);
	signal p153_out : STD_LOGIC;
	signal p154_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p154_out : STD_LOGIC;
	signal p155_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p155_out : STD_LOGIC;
	signal p156_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p156_out : STD_LOGIC;
	signal p157_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p157_out : STD_LOGIC;
	signal p158_in : STD_LOGIC_VECTOR(0 to 51 - 1);
	signal p158_out : STD_LOGIC;
	signal p159_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p159_out : STD_LOGIC;
	signal p160_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p160_out : STD_LOGIC;
	signal p161_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p161_out : STD_LOGIC;
	signal p162_in : STD_LOGIC_VECTOR(0 to 54 - 1);
	signal p162_out : STD_LOGIC;
	signal p163_in : STD_LOGIC_VECTOR(0 to 59 - 1);
	signal p163_out : STD_LOGIC;
	signal p164_in : STD_LOGIC_VECTOR(0 to 54 - 1);
	signal p164_out : STD_LOGIC;
	signal p165_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p165_out : STD_LOGIC;
	signal p166_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p166_out : STD_LOGIC;
	signal p167_in : STD_LOGIC_VECTOR(0 to 47 - 1);
	signal p167_out : STD_LOGIC;
	signal p168_in : STD_LOGIC_VECTOR(0 to 51 - 1);
	signal p168_out : STD_LOGIC;
	signal p169_in : STD_LOGIC_VECTOR(0 to 44 - 1);
	signal p169_out : STD_LOGIC;
	signal p170_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p170_out : STD_LOGIC;
	signal p171_in : STD_LOGIC_VECTOR(0 to 63 - 1);
	signal p171_out : STD_LOGIC;
	signal p172_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p172_out : STD_LOGIC;
	signal p173_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p173_out : STD_LOGIC;
	signal p174_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p174_out : STD_LOGIC;
	signal p175_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p175_out : STD_LOGIC;
	signal p176_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p176_out : STD_LOGIC;
	signal p177_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p177_out : STD_LOGIC;
	signal p178_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p178_out : STD_LOGIC;
	signal p179_in : STD_LOGIC_VECTOR(0 to 81 - 1);
	signal p179_out : STD_LOGIC;
	signal p180_in : STD_LOGIC_VECTOR(0 to 75 - 1);
	signal p180_out : STD_LOGIC;
	signal p181_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p181_out : STD_LOGIC;
	signal p182_in : STD_LOGIC_VECTOR(0 to 50 - 1);
	signal p182_out : STD_LOGIC;
	signal p183_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p183_out : STD_LOGIC;
	signal p184_in : STD_LOGIC_VECTOR(0 to 46 - 1);
	signal p184_out : STD_LOGIC;
	signal p185_in : STD_LOGIC_VECTOR(0 to 56 - 1);
	signal p185_out : STD_LOGIC;
	signal p186_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p186_out : STD_LOGIC;
	signal p187_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p187_out : STD_LOGIC;
	signal p188_in : STD_LOGIC_VECTOR(0 to 50 - 1);
	signal p188_out : STD_LOGIC;
	signal p189_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p189_out : STD_LOGIC;
	signal p190_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p190_out : STD_LOGIC;
	signal p191_in : STD_LOGIC_VECTOR(0 to 54 - 1);
	signal p191_out : STD_LOGIC;
	signal p192_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p192_out : STD_LOGIC;
	signal p193_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p193_out : STD_LOGIC;
	signal p194_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p194_out : STD_LOGIC;
	signal p195_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p195_out : STD_LOGIC;
	signal p196_in : STD_LOGIC_VECTOR(0 to 63 - 1);
	signal p196_out : STD_LOGIC;
	signal p197_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p197_out : STD_LOGIC;
	signal p198_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p198_out : STD_LOGIC;
	signal p199_in : STD_LOGIC_VECTOR(0 to 47 - 1);
	signal p199_out : STD_LOGIC;
	signal p200_in : STD_LOGIC_VECTOR(0 to 48 - 1);
	signal p200_out : STD_LOGIC;
	signal p201_in : STD_LOGIC_VECTOR(0 to 48 - 1);
	signal p201_out : STD_LOGIC;
	signal p202_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p202_out : STD_LOGIC;
	signal p203_in : STD_LOGIC_VECTOR(0 to 50 - 1);
	signal p203_out : STD_LOGIC;
	signal p204_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p204_out : STD_LOGIC;
	signal p205_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p205_out : STD_LOGIC;
	signal p206_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p206_out : STD_LOGIC;
	signal p207_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p207_out : STD_LOGIC;
	signal p208_in : STD_LOGIC_VECTOR(0 to 86 - 1);
	signal p208_out : STD_LOGIC;
	signal p209_in : STD_LOGIC_VECTOR(0 to 45 - 1);
	signal p209_out : STD_LOGIC;
	signal p210_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p210_out : STD_LOGIC;
	signal p211_in : STD_LOGIC_VECTOR(0 to 62 - 1);
	signal p211_out : STD_LOGIC;
	signal p212_in : STD_LOGIC_VECTOR(0 to 46 - 1);
	signal p212_out : STD_LOGIC;
	signal p213_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p213_out : STD_LOGIC;
	signal p214_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p214_out : STD_LOGIC;
	signal p215_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p215_out : STD_LOGIC;
	signal p216_in : STD_LOGIC_VECTOR(0 to 58 - 1);
	signal p216_out : STD_LOGIC;
	signal p217_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p217_out : STD_LOGIC;
	signal p218_in : STD_LOGIC_VECTOR(0 to 60 - 1);
	signal p218_out : STD_LOGIC;
	signal p219_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p219_out : STD_LOGIC;
	signal p220_in : STD_LOGIC_VECTOR(0 to 75 - 1);
	signal p220_out : STD_LOGIC;
	signal p221_in : STD_LOGIC_VECTOR(0 to 48 - 1);
	signal p221_out : STD_LOGIC;
	signal p222_in : STD_LOGIC_VECTOR(0 to 72 - 1);
	signal p222_out : STD_LOGIC;
	signal p223_in : STD_LOGIC_VECTOR(0 to 64 - 1);
	signal p223_out : STD_LOGIC;
	signal p224_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p224_out : STD_LOGIC;
	signal p225_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p225_out : STD_LOGIC;
	signal p226_in : STD_LOGIC_VECTOR(0 to 49 - 1);
	signal p226_out : STD_LOGIC;
	signal p227_in : STD_LOGIC_VECTOR(0 to 58 - 1);
	signal p227_out : STD_LOGIC;
	signal p228_in : STD_LOGIC_VECTOR(0 to 46 - 1);
	signal p228_out : STD_LOGIC;
	signal p229_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p229_out : STD_LOGIC;
	signal p230_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p230_out : STD_LOGIC;
	signal p231_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p231_out : STD_LOGIC;
	signal p232_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p232_out : STD_LOGIC;
	signal p233_in : STD_LOGIC_VECTOR(0 to 67 - 1);
	signal p233_out : STD_LOGIC;
	signal p234_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p234_out : STD_LOGIC;
	signal p235_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p235_out : STD_LOGIC;
	signal p236_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p236_out : STD_LOGIC;
	signal p237_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p237_out : STD_LOGIC;
	signal p238_in : STD_LOGIC_VECTOR(0 to 50 - 1);
	signal p238_out : STD_LOGIC;
	signal p239_in : STD_LOGIC_VECTOR(0 to 60 - 1);
	signal p239_out : STD_LOGIC;
	signal p240_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p240_out : STD_LOGIC;
	signal p241_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p241_out : STD_LOGIC;
	signal p242_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p242_out : STD_LOGIC;
	signal p243_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p243_out : STD_LOGIC;
	signal p244_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p244_out : STD_LOGIC;
	signal p245_in : STD_LOGIC_VECTOR(0 to 74 - 1);
	signal p245_out : STD_LOGIC;
	signal p246_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p246_out : STD_LOGIC;
	signal p247_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p247_out : STD_LOGIC;
	signal p248_in : STD_LOGIC_VECTOR(0 to 64 - 1);
	signal p248_out : STD_LOGIC;
	signal p249_in : STD_LOGIC_VECTOR(0 to 67 - 1);
	signal p249_out : STD_LOGIC;
	signal p250_in : STD_LOGIC_VECTOR(0 to 75 - 1);
	signal p250_out : STD_LOGIC;
	signal p251_in : STD_LOGIC_VECTOR(0 to 44 - 1);
	signal p251_out : STD_LOGIC;
	signal p252_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p252_out : STD_LOGIC;
	signal p253_in : STD_LOGIC_VECTOR(0 to 66 - 1);
	signal p253_out : STD_LOGIC;
	signal p254_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p254_out : STD_LOGIC;
	signal p255_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p255_out : STD_LOGIC;
	
    
    -- Dummies
    signal dummy0 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy1 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy2 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy3 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy4 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy5 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy6 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy7 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy8 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy9 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy10 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy11 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy12 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy13 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy14 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy15 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy16 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy17 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy18 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy19 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy20 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy21 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy22 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy23 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy24 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy25 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy26 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy27 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy28 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy29 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy30 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy31 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy32 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy33 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy34 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy35 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy36 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy37 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy38 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy39 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy40 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy41 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy42 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy43 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy44 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy45 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy46 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy47 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy48 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy49 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy50 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy51 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy52 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy53 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy54 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy55 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy56 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy57 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy58 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy59 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy60 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy61 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy62 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy63 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy64 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy65 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy66 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy67 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy68 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy69 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy70 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy71 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy72 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy73 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy74 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy75 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy76 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy77 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy78 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy79 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy80 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy81 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy82 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy83 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy84 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy85 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy86 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy87 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy88 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy89 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy90 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy91 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy92 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy93 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy94 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy95 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy96 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy97 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy98 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy99 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy100 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy101 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy102 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy103 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy104 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy105 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy106 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy107 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy108 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy109 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy110 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy111 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy112 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy113 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy114 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy115 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy116 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy117 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy118 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy119 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy120 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy121 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy122 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy123 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy124 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy125 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy126 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy127 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy128 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy129 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy130 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy131 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy132 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy133 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy134 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy135 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy136 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy137 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy138 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy139 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy140 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy141 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy142 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy143 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy144 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy145 : STD_LOGIC_VECTOR(0 to 12 - 2);
	signal dummy146 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy147 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy148 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy149 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy150 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy151 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy152 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy153 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy154 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy155 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy156 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy157 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy158 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy159 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy160 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy161 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy162 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy163 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy164 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy165 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy166 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy167 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy168 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy169 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy170 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy171 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy172 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy173 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy174 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy175 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy176 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy177 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy178 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy179 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy180 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy181 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy182 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy183 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy184 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy185 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy186 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy187 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy188 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy189 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy190 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy191 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy192 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy193 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy194 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy195 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy196 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy197 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy198 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy199 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy200 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy201 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy202 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy203 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy204 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy205 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy206 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy207 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy208 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy209 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy210 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy211 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy212 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy213 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy214 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy215 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy216 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy217 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy218 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy219 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy220 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy221 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy222 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy223 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy224 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy225 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy226 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy227 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy228 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy229 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy230 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy231 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy232 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy233 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy234 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy235 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy236 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy237 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy238 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy239 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy240 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy241 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy242 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy243 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy244 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy245 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy246 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy247 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy248 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy249 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy250 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy251 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy252 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy253 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy254 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy255 : STD_LOGIC_VECTOR(0 to 13 - 2);
	 

begin

    
    p0_in <= x(249) & x(276) & x(277) & x(294) & x(304) & x(305) & x(306) & x(330) & x(331) & x(333) & x(334) & x(338) & x(357) & x(358) & x(359) & x(360) & x(362) & x(366) & x(370) & x(386) & x(387) & x(388) & x(390) & x(397) & x(418) & x(424) & x(446) & x(474) & x(501) & x(529) & x(707) & x(708) & x(709) & x(739) & x(742) & x(743) & x(744) & x(745) & x(746);
    y(0) <= not(p0_out);
    p0 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111100111000011000010101111111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 3,
            B => 119,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p0_in,
            y(0) => p0_out,
            y(1 to 14 - 1) => dummy0
        );


    p1_in <= x(178) & x(192) & x(198) & x(220) & x(228) & x(242) & x(248) & x(249) & x(270) & x(276) & x(277) & x(297) & x(298) & x(299) & x(300) & x(304) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(333) & x(334) & x(342) & x(351) & x(357) & x(358) & x(359) & x(360) & x(362) & x(369) & x(370) & x(371) & x(378) & x(379) & x(386) & x(387) & x(388) & x(390) & x(397) & x(405) & x(406) & x(407) & x(415) & x(416) & x(418) & x(425) & x(433) & x(442) & x(443) & x(450) & x(584) & x(611) & x(666) & x(682) & x(692) & x(696) & x(717);
    y(1) <= not(p1_out);
    p1 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10001100100111100011110010111101110011101000110101110001000",
            TABLE => "01110001000100000001000000000000111101110111000101110001000100000111000100011000000110001000111011100111011100010111000100011000011010011001011010010110011010011001011001101001011010011001011011010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100100000000100000001000000011101000100000001110100011101000111111100001011110000001100000011110100010000001111010001110100001111110011010011001011010010110011010011001011001101001011010011001011000000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100100000001000101110000000000000001000101110111111100000001000101111000000100010111111010001000000100010111011111101000000100010111011010011001011010010110011010011001011001101001011010011001011000001000100011101000111011101111000000000000100000001000100011100001100010001110100011101110011101110001000110000001100010001110011010011001011010010110011010011001011001101001011010011001011000000000001000000010000010110010001000001011001010110010111110110100110100100100001001001011001000100100101100101011001011011011100101100110100101101001100101100110100110010110100101100110100101001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011000001000100011101000111011101111000000000000100000001000100011100001100010001110100011101110011101110001000110000001100010001110011010011001011010010110011010011001011001101001011010011001011011101000111111101000000011101000111010000111111010000001111010000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 1,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p1_in,
            y(0) => p1_out,
            y(1 to 13 - 1) => dummy1
        );


    p2_in <= x(192) & x(220) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(310) & x(321) & x(322) & x(333) & x(334) & x(357) & x(426) & x(454) & x(486) & x(666) & x(697) & x(707);
    y(2) <= not(p2_out);
    p2 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000000001111110",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 3,
            B => -133,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p2_in,
            y(0) => p2_out,
            y(1 to 13 - 1) => dummy2
        );


    p3_in <= x(63) & x(106) & x(260) & x(294) & x(295) & x(313) & x(314) & x(315) & x(341) & x(342) & x(369) & x(370) & x(502);
    y(3) <= not(p3_out);
    p3 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001100000001",
            TABLE => "1011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => -68,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p3_in,
            y(0) => p3_out,
            y(1 to 12 - 1) => dummy3
        );


    p4_in <= x(40) & x(162) & x(183) & x(276) & x(304) & x(339) & x(342) & x(355) & x(366) & x(367) & x(369) & x(381) & x(382) & x(403) & x(404) & x(409) & x(410) & x(436) & x(665) & x(679) & x(692) & x(707);
    y(4) <= not(p4_out);
    p4 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101111011100000000101",
            TABLE => "0000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010100110100000100010011010010010001101001100101100000000000000000",
            SHIFT => 3,
            B => 52,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p4_in,
            y(0) => p4_out,
            y(1 to 13 - 1) => dummy4
        );


    p5_in <= x(157) & x(190) & x(191) & x(205) & x(211) & x(218) & x(233) & x(243) & x(248) & x(276) & x(277) & x(294) & x(305) & x(322) & x(328) & x(330) & x(331) & x(332) & x(350) & x(358) & x(359) & x(360) & x(375) & x(378) & x(379) & x(399) & x(400) & x(401) & x(402) & x(407) & x(418) & x(428) & x(446) & x(466) & x(467) & x(473) & x(494) & x(515) & x(528) & x(604) & x(607) & x(611) & x(635) & x(664) & x(665) & x(695) & x(697) & x(707) & x(718) & x(719) & x(720) & x(721) & x(735) & x(739) & x(740) & x(741) & x(742) & x(745) & x(746);
    y(5) <= not(p5_out);
    p5 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11110111111010000000001001111011111110111111101000000000000",
            TABLE => "00000000000001000000010001001101000001000100110101001101110111111011001000100100001001000100110100100100010011010100110111011011011010011001011010010110011010011001011001101001011010011001011000000000000000100000001000101011000000100010101100101011101111111101010001000010010000100010101101000010001010110010101110111101011010011001011010010110011010011001011001101001011010011001011011101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011011111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011000000010001010110010101110111111000000000000001000000010001010110100001000101011001010111011110111010100010000100100001000101011100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000001000101110000000000000001000101110111111100000001000101111000000100010111111010001000000100010111011111101000000100010111011010011001011010010110011010011001011001101001011010011001011000000000001000000010000010110010001000001011001010110010111110110100110100100100001001001011001000100100101100101011001011011011100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 2,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p5_in,
            y(0) => p5_out,
            y(1 to 14 - 1) => dummy5
        );


    p6_in <= x(89) & x(98) & x(99) & x(117) & x(118) & x(121) & x(122) & x(133) & x(134) & x(135) & x(147) & x(152) & x(153) & x(163) & x(180) & x(181) & x(182) & x(191) & x(192) & x(219) & x(220) & x(247) & x(248) & x(275) & x(276) & x(277) & x(317) & x(344) & x(350) & x(369) & x(371) & x(390) & x(391) & x(443) & x(474) & x(475) & x(502) & x(522) & x(564) & x(592) & x(619) & x(668) & x(720) & x(721);
    y(6) <= not(p6_out);
    p6 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111110001110111000000000001001101111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 2,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p6_in,
            y(0) => p6_out,
            y(1 to 13 - 1) => dummy6
        );


    p7_in <= x(64) & x(66) & x(136) & x(144) & x(145) & x(171) & x(174) & x(184) & x(188) & x(199) & x(200) & x(201) & x(212) & x(228) & x(248) & x(256) & x(276) & x(277) & x(283) & x(295) & x(296) & x(297) & x(304) & x(305) & x(306) & x(310) & x(311) & x(316) & x(324) & x(325) & x(333) & x(334) & x(338) & x(339) & x(352) & x(366) & x(411) & x(439) & x(474) & x(475) & x(542) & x(582) & x(583) & x(610) & x(666) & x(667) & x(676) & x(695) & x(705) & x(708) & x(723) & x(724) & x(774);
    y(7) <= not(p7_out);
    p7 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00011110011101010011110001101100111111110000001011001",
            TABLE => "01111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011000010111000000010000000100000000011111110001011100010111000000010001011110000001100000011110100001111110000101110001011110000001100101100110100101101001100101100110100110010110100101100110100110001110000010001110111110001110000010000000000010001110000010001000111000011000111001111000111000011000011100011000111000011000100101100110100101101001100101100110100110010110100101100110100100000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100100010000011100010111000111110111000000000001000000010000011100010001100001110001011100011110011110001110000110000001100001110001100101100110100101101001100101100110100110010110100101100110100100010111011111110000000100010111000000010001011100000000000000010001011101111110100000010001011110000001000101111110100010000001100101100110100101101001100101100110100110010110100101100110100100000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100111111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011001000000110101001101010011111101010000101101010011010100101111010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 3,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p7_in,
            y(0) => p7_out,
            y(1 to 14 - 1) => dummy7
        );


    p8_in <= x(65) & x(66) & x(93) & x(94) & x(198) & x(239) & x(240) & x(267) & x(268) & x(338) & x(473) & x(501) & x(528) & x(529) & x(605) & x(631) & x(634) & x(658) & x(659) & x(660) & x(705);
    y(8) <= not(p8_out);
    p8 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000001111000000000001",
            TABLE => "111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001110101001001011011111111",
            SHIFT => 3,
            B => -77,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p8_in,
            y(0) => p8_out,
            y(1 to 13 - 1) => dummy8
        );


    p9_in <= x(68) & x(78) & x(192) & x(198) & x(220) & x(248) & x(249) & x(257) & x(276) & x(277) & x(302) & x(304) & x(305) & x(306) & x(322) & x(329) & x(330) & x(331) & x(350) & x(358) & x(361) & x(389) & x(390) & x(418) & x(446) & x(453) & x(454) & x(474) & x(475) & x(502) & x(531) & x(675) & x(697) & x(719);
    y(9) <= not(p9_out);
    p9 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001000100100001110111111111111010",
            TABLE => "1110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101101011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010010000010110010001001001011001001101001100101100000000000000000",
            SHIFT => 3,
            B => 21,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p9_in,
            y(0) => p9_out,
            y(1 to 14 - 1) => dummy9
        );


    p10_in <= x(135) & x(163) & x(262) & x(263) & x(289) & x(290) & x(309) & x(310) & x(315) & x(332) & x(338) & x(344) & x(366) & x(412) & x(433) & x(434) & x(435) & x(440) & x(459) & x(460) & x(461) & x(473) & x(501) & x(529) & x(611) & x(688);
    y(10) <= not(p10_out);
    p10 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000010000111011100001",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 2,
            B => -53,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p10_in,
            y(0) => p10_out,
            y(1 to 12 - 1) => dummy10
        );


    p11_in <= x(171) & x(183) & x(200) & x(228) & x(267) & x(276) & x(294) & x(295) & x(310) & x(311) & x(316) & x(339) & x(342) & x(358) & x(359) & x(386) & x(387) & x(389) & x(418) & x(446) & x(474) & x(502) & x(691) & x(772) & x(773) & x(774);
    y(11) <= not(p11_out);
    p11 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01000100001011111000001000",
            TABLE => "110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 3,
            B => -65,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p11_in,
            y(0) => p11_out,
            y(1 to 13 - 1) => dummy11
        );


    p12_in <= x(66) & x(71) & x(72) & x(136) & x(165) & x(192) & x(220) & x(248) & x(249) & x(276) & x(277) & x(289) & x(305) & x(306) & x(311) & x(315) & x(316) & x(329) & x(330) & x(331) & x(333) & x(334) & x(341) & x(350) & x(351) & x(359) & x(360) & x(379) & x(387) & x(388) & x(401) & x(406) & x(407) & x(416) & x(424) & x(425) & x(426) & x(427) & x(428) & x(453) & x(454) & x(455) & x(481) & x(482) & x(501) & x(511) & x(557) & x(687) & x(690) & x(691) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(724) & x(748) & x(750);
    y(12) <= not(p12_out);
    p12 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000100111000001101110011111111111111000000000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 2,
            B => -50,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p12_in,
            y(0) => p12_out,
            y(1 to 14 - 1) => dummy12
        );


    p13_in <= x(145) & x(247) & x(266) & x(276) & x(293) & x(294) & x(295) & x(304) & x(305) & x(321) & x(327) & x(418) & x(435) & x(473) & x(474) & x(501) & x(502) & x(507) & x(528) & x(557) & x(583) & x(584) & x(610) & x(611) & x(613) & x(638) & x(675) & x(697) & x(706);
    y(13) <= not(p13_out);
    p13 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000000001010000100000000101",
            TABLE => "11101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011011111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011011010100010000000100000000000000111111011101010011010100010000001101010001000010010000100010101110111101110101001101010001000010100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111011111010011010100110100000100110110110100110101001101001001001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -137,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p13_in,
            y(0) => p13_out,
            y(1 to 14 - 1) => dummy13
        );


    p14_in <= x(192) & x(193) & x(221) & x(248) & x(249) & x(276) & x(277) & x(305) & x(330) & x(331) & x(347) & x(377) & x(390) & x(418) & x(446) & x(474) & x(486) & x(502) & x(514) & x(517) & x(528) & x(529) & x(557) & x(675) & x(676) & x(694) & x(695) & x(705) & x(706) & x(707) & x(708) & x(709) & x(722) & x(723) & x(732) & x(733);
    y(14) <= not(p14_out);
    p14 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111110011000000000001111111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 108,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p14_in,
            y(0) => p14_out,
            y(1 to 15 - 1) => dummy14
        );


    p15_in <= x(66) & x(95) & x(192) & x(220) & x(221) & x(248) & x(249) & x(276) & x(277) & x(295) & x(305) & x(330) & x(331) & x(332) & x(357) & x(358) & x(359) & x(360) & x(366) & x(386) & x(387) & x(388) & x(416) & x(514);
    y(15) <= not(p15_out);
    p15 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110000000001111111011111",
            TABLE => "100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => 23,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p15_in,
            y(0) => p15_out,
            y(1 to 13 - 1) => dummy15
        );


    p16_in <= x(92) & x(204) & x(210) & x(220) & x(248) & x(249) & x(260) & x(276) & x(277) & x(278) & x(284) & x(305) & x(306) & x(339) & x(350) & x(351) & x(378) & x(379) & x(389) & x(685) & x(695);
    y(16) <= not(p16_out);
    p16 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001000000000001111001",
            TABLE => "111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001110101001001011011111111",
            SHIFT => 3,
            B => -106,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p16_in,
            y(0) => p16_out,
            y(1 to 13 - 1) => dummy16
        );


    p17_in <= x(93) & x(95) & x(96) & x(108) & x(118) & x(153) & x(163) & x(191) & x(192) & x(219) & x(220) & x(221) & x(238) & x(248) & x(249) & x(266) & x(267) & x(276) & x(277) & x(304) & x(305) & x(306) & x(316) & x(317) & x(318) & x(327) & x(328) & x(329) & x(330) & x(331) & x(333) & x(334) & x(342) & x(343) & x(344) & x(345) & x(346) & x(347) & x(357) & x(358) & x(359) & x(360) & x(370) & x(389) & x(418) & x(453) & x(454) & x(474) & x(475) & x(502) & x(549) & x(613) & x(661) & x(668) & x(705) & x(720) & x(734) & x(736) & x(737) & x(738) & x(741) & x(742) & x(745) & x(746) & x(747);
    y(17) <= not(p17_out);
    p17 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111100000010011000000001111100000000111101111111110111111111111",
            TABLE => "00000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100101011000000100000001000000000101111110010101100101011000000100010101101000010010000101101010010111101001010110010101101000010011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100000001000101110001011101111111000000000000000100000001000101111000000100010111000101110111111011101000100000011000000100010111011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100010111011111110000000100010111000000010001011100000000000000010001011101111110100000010001011110000001000101111110100010000001100101100110100101101001100101100110100110010110100101100110100100000001000101110001011101111111000000000000000100000001000101111000000100010111000101110111111011101000100000011000000100010111011010011001011010010110011010011001011001101001011010011001011000000000000001000000010001001101000001000100110101001101110111111011001000100100001001000100110100100100010011010100110111011011011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000001000101110001011101111111100000010001011100010111011111100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 2,
            B => 45,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p17_in,
            y(0) => p17_out,
            y(1 to 14 - 1) => dummy17
        );


    p18_in <= x(179) & x(206) & x(248) & x(276) & x(277) & x(294) & x(295) & x(305) & x(322) & x(357) & x(358) & x(359) & x(360) & x(387) & x(389) & x(494) & x(522) & x(654) & x(657) & x(685) & x(686) & x(742) & x(745) & x(746);
    y(18) <= not(p18_out);
    p18 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110000000111111111111000",
            TABLE => "100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p18_in,
            y(0) => p18_out,
            y(1 to 13 - 1) => dummy18
        );


    p19_in <= x(152) & x(267) & x(268) & x(269) & x(295) & x(296) & x(310) & x(338) & x(342) & x(359) & x(366) & x(370) & x(371) & x(398) & x(418) & x(446) & x(473) & x(474) & x(501) & x(502) & x(508) & x(528) & x(529) & x(557) & x(697) & x(742);
    y(19) <= not(p19_out);
    p19 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000000110111000000000000",
            TABLE => "111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 3,
            B => -71,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p19_in,
            y(0) => p19_out,
            y(1 to 13 - 1) => dummy19
        );


    p20_in <= x(35) & x(50) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(79) & x(89) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(101) & x(102) & x(104) & x(107) & x(108) & x(192) & x(219) & x(220) & x(228) & x(247) & x(248) & x(249) & x(275) & x(276) & x(277) & x(304) & x(305) & x(306) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(334) & x(354) & x(359) & x(360) & x(361) & x(370) & x(388) & x(396) & x(397) & x(445) & x(473) & x(474) & x(529) & x(609) & x(611) & x(636) & x(638) & x(665) & x(666) & x(679) & x(692) & x(739) & x(745);
    y(20) <= not(p20_out);
    p20 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000000000000000000000001110111111111000000010000101100001111110100",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101101111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101101000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011000111000001000100011100001100010010110011010010000000000000000",
            SHIFT => 3,
            B => -122,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p20_in,
            y(0) => p20_out,
            y(1 to 15 - 1) => dummy20
        );


    p21_in <= x(41) & x(98) & x(99) & x(101) & x(108) & x(136) & x(152) & x(160) & x(161) & x(162) & x(163) & x(181) & x(192) & x(210) & x(220) & x(221) & x(247) & x(248) & x(249) & x(276) & x(277) & x(299) & x(300) & x(302) & x(305) & x(306) & x(323) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(333) & x(334) & x(358) & x(359) & x(360) & x(379) & x(387) & x(388) & x(406) & x(415) & x(416) & x(418) & x(434) & x(443) & x(461) & x(489) & x(517) & x(593) & x(611) & x(676) & x(705) & x(706);
    y(21) <= not(p21_out);
    p21 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000010111101011111110001110000001100010010011011101000",
            TABLE => "1111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010010000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101101011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010010100110111011111000001000100110100000100010011010000000000000100010011011101101100100100010011010010010001001101101100100010010001101001100101101001011001101001100101100110100101101001100101100000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 2,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p21_in,
            y(0) => p21_out,
            y(1 to 13 - 1) => dummy21
        );


    p22_in <= x(215) & x(228) & x(247) & x(276) & x(304) & x(320) & x(343) & x(348) & x(351) & x(352) & x(370) & x(380) & x(390) & x(418) & x(446) & x(474) & x(507) & x(528) & x(529) & x(535) & x(557) & x(611) & x(622);
    y(22) <= not(p22_out);
    p22 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10111000000011110110111",
            TABLE => "00000010001010110000000000000010001010111011111100000010001010110100001000101011110101000100001000101011101111010100001000101011100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100000000000001000000010001001101000001000100110101001101110111111011001000100100001001000100110100100100010011010100110111011011011010011001011010010110011010011001011001101001011010011001011000010111000000010111111100010111000101111000000101111110000101111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => 62,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p22_in,
            y(0) => p22_out,
            y(1 to 13 - 1) => dummy22
        );


    p23_in <= x(117) & x(145) & x(147) & x(161) & x(219) & x(228) & x(247) & x(248) & x(276) & x(294) & x(314) & x(315) & x(321) & x(322) & x(338) & x(341) & x(342) & x(352) & x(366) & x(375) & x(377) & x(380) & x(381) & x(382) & x(403) & x(404) & x(409) & x(410) & x(436) & x(460) & x(464) & x(507) & x(535) & x(660) & x(693) & x(694) & x(739);
    y(23) <= not(p23_out);
    p23 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001101111111111101000000000000001001",
            TABLE => "1011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 2,
            B => 19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p23_in,
            y(0) => p23_out,
            y(1 to 13 - 1) => dummy23
        );


    p24_in <= x(35) & x(40) & x(41) & x(46) & x(50) & x(78) & x(95) & x(107) & x(108) & x(116) & x(162) & x(190) & x(192) & x(218) & x(220) & x(221) & x(243) & x(246) & x(247) & x(248) & x(249) & x(263) & x(275) & x(276) & x(277) & x(304) & x(305) & x(306) & x(326) & x(327) & x(328) & x(329) & x(330) & x(331) & x(333) & x(334) & x(338) & x(339) & x(353) & x(357) & x(358) & x(359) & x(360) & x(362) & x(366) & x(387) & x(388) & x(390) & x(412) & x(418) & x(451) & x(486) & x(508) & x(509) & x(510) & x(513) & x(514) & x(515) & x(538) & x(584) & x(611) & x(666) & x(688) & x(697) & x(712);
    y(24) <= not(p24_out);
    p24 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000001111111111111111110000001111000001100111101110001111011",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100111110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100110000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100101000000110101001101010011111101000000000100000001000000110101000100001011010100110101001011110100101011010000100100001011010100011010011001011010010110011010011001011001101001011010011001011000000000000100000001000001110001000100000111000101110001111101111000111000011000000110000111000100011000011100010111000111100111011010011001011010010110011010011001011001101001011010011001011001110001000100000001000000000000111101110111000101110001000100000111000100011000000110001000111011100111011100010111000100011000011010011001011010010110011010011001011001101001011010011001011000010000011100010111000111110111000110000111000101110001111001111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 2,
            B => 69,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p24_in,
            y(0) => p24_out,
            y(1 to 14 - 1) => dummy24
        );


    p25_in <= x(228) & x(238) & x(249) & x(256) & x(277) & x(283) & x(305) & x(310) & x(311) & x(312) & x(323) & x(324) & x(338) & x(339) & x(358) & x(359) & x(360) & x(368) & x(403) & x(410) & x(422) & x(445) & x(464) & x(473) & x(474) & x(485) & x(487) & x(500) & x(501) & x(514) & x(527) & x(528) & x(542) & x(600) & x(601) & x(628) & x(677) & x(678);
    y(25) <= not(p25_out);
    p25 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10111111111111000101101000000000000011",
            TABLE => "000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 3,
            B => 39,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p25_in,
            y(0) => p25_out,
            y(1 to 14 - 1) => dummy25
        );


    p26_in <= x(136) & x(192) & x(220) & x(248) & x(249) & x(266) & x(276) & x(277) & x(305) & x(306) & x(329) & x(330) & x(331) & x(332) & x(334) & x(358) & x(359) & x(360) & x(386) & x(387) & x(388) & x(389) & x(391) & x(418) & x(473) & x(474) & x(501) & x(528) & x(529) & x(557) & x(697);
    y(26) <= not(p26_out);
    p26 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000010000111101111111111111111",
            TABLE => "1111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101101111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => 66,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p26_in,
            y(0) => p26_out,
            y(1 to 14 - 1) => dummy26
        );


    p27_in <= x(160) & x(161) & x(162) & x(163) & x(276) & x(277) & x(295) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(333) & x(338) & x(339) & x(358) & x(359) & x(360) & x(366) & x(386) & x(387) & x(388) & x(391) & x(418) & x(536) & x(696) & x(724) & x(750);
    y(27) <= not(p27_out);
    p27 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000011110001110111000000",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100101111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011001110001000100000001000000000000111101110111000101110001000100000111000100011000000110001000111011100111011100010111000100011000011010011001011010010110011010011001011001101001011010011001011000000010001010110000000000000010001010111011111100000010001010110100001000101011110101000100001000101011101111010100001000101011100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -84,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p27_in,
            y(0) => p27_out,
            y(1 to 14 - 1) => dummy27
        );


    p28_in <= x(65) & x(66) & x(91) & x(93) & x(108) & x(136) & x(191) & x(192) & x(198) & x(220) & x(221) & x(248) & x(249) & x(276) & x(277) & x(305) & x(306) & x(329) & x(330) & x(331) & x(332) & x(334) & x(343) & x(346) & x(347) & x(348) & x(357) & x(358) & x(359) & x(360) & x(370) & x(371) & x(387) & x(388) & x(396) & x(418) & x(454) & x(473) & x(474) & x(501) & x(514) & x(515) & x(675);
    y(28) <= not(p28_out);
    p28 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000011101111111100001111100001100100000001",
            TABLE => "1111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101101000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p28_in,
            y(0) => p28_out,
            y(1 to 14 - 1) => dummy28
        );


    p29_in <= x(91) & x(93) & x(94) & x(95) & x(108) & x(192) & x(248) & x(249) & x(276) & x(277) & x(305) & x(322) & x(329) & x(330) & x(333) & x(338) & x(342) & x(343) & x(344) & x(345) & x(348) & x(349) & x(350) & x(351) & x(360) & x(369) & x(370) & x(371) & x(372) & x(376) & x(377) & x(378) & x(389) & x(391) & x(396) & x(417) & x(418) & x(473) & x(474) & x(486) & x(487) & x(500) & x(501) & x(514) & x(515) & x(516) & x(528) & x(529) & x(542) & x(666) & x(697) & x(717) & x(738) & x(739) & x(740) & x(741) & x(742) & x(744) & x(745) & x(746) & x(747) & x(770) & x(774);
    y(29) <= not(p29_out);
    p29 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111110000000110100000000100000001101111111111111111111111111111",
            TABLE => "000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 2,
            B => 66,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p29_in,
            y(0) => p29_out,
            y(1 to 14 - 1) => dummy29
        );


    p30_in <= x(292) & x(305) & x(333) & x(354) & x(358) & x(380) & x(415) & x(416) & x(435) & x(444) & x(453) & x(463) & x(656) & x(657) & x(658);
    y(30) <= not(p30_out);
    p30 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011101001001111",
            TABLE => "000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 3,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p30_in,
            y(0) => p30_out,
            y(1 to 13 - 1) => dummy30
        );


    p31_in <= x(64) & x(66) & x(136) & x(163) & x(164) & x(171) & x(172) & x(183) & x(192) & x(193) & x(194) & x(201) & x(220) & x(221) & x(222) & x(242) & x(243) & x(244) & x(245) & x(248) & x(249) & x(276) & x(277) & x(304) & x(305) & x(306) & x(311) & x(320) & x(328) & x(329) & x(330) & x(331) & x(332) & x(339) & x(343) & x(346) & x(347) & x(356) & x(357) & x(358) & x(359) & x(360) & x(366) & x(368) & x(370) & x(371) & x(387) & x(388) & x(389) & x(396) & x(405) & x(406) & x(407) & x(422) & x(433) & x(434) & x(435) & x(439) & x(440) & x(442) & x(443) & x(467) & x(468) & x(494) & x(495) & x(496) & x(497) & x(514) & x(515) & x(535) & x(602) & x(648) & x(649) & x(675) & x(676) & x(677) & x(679) & x(690) & x(704) & x(705) & x(706) & x(707) & x(708) & x(709) & x(710);
    y(31) <= not(p31_out);
    p31 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100000100000000000000000000111110000111110000111011101110000000000110100000010000000",
            TABLE => "1000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101101111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101101111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 2,
            B => -127,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p31_in,
            y(0) => p31_out,
            y(1 to 14 - 1) => dummy31
        );


    p32_in <= x(35) & x(62) & x(63) & x(65) & x(66) & x(68) & x(91) & x(135) & x(144) & x(145) & x(162) & x(192) & x(221) & x(228) & x(248) & x(249) & x(276) & x(277) & x(287) & x(289) & x(305) & x(306) & x(329) & x(330) & x(331) & x(332) & x(357) & x(358) & x(359) & x(360) & x(361) & x(485) & x(501) & x(528) & x(529) & x(571) & x(584) & x(598) & x(599) & x(600) & x(649);
    y(32) <= not(p32_out);
    p32 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000110001000000001111111111000000000",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100110001110111011110000100010001110000010001000111000000000000010001000111011100111000110001000111000011000100011100111000100011000100101100110100101101001100101100110100110010110100101100110100111101000100000001111111011101000100000000000000011101000100000001110100010000001011111101110100010000001000101111110100010000001011010011001011010010110011010011001011001101001011010011001011011110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100110000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -109,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p32_in,
            y(0) => p32_out,
            y(1 to 14 - 1) => dummy32
        );


    p33_in <= x(35) & x(40) & x(41) & x(63) & x(64) & x(134) & x(135) & x(155) & x(156) & x(208) & x(230) & x(257) & x(276) & x(342) & x(361) & x(362) & x(368) & x(369) & x(370) & x(389) & x(390) & x(418) & x(446) & x(463) & x(474) & x(475) & x(492) & x(502) & x(544) & x(636) & x(662) & x(663) & x(695) & x(705) & x(722) & x(723) & x(742);
    y(33) <= not(p33_out);
    p33 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111111001001100111000000000100011111",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => 21,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p33_in,
            y(0) => p33_out,
            y(1 to 14 - 1) => dummy33
        );


    p34_in <= x(44) & x(116) & x(158) & x(189) & x(190) & x(217) & x(260) & x(263) & x(276) & x(287) & x(290) & x(291) & x(292) & x(310) & x(338) & x(339) & x(362) & x(366) & x(377) & x(390) & x(418) & x(446) & x(474) & x(656) & x(658) & x(659) & x(660) & x(686) & x(694) & x(695) & x(732) & x(733) & x(774);
    y(34) <= not(p34_out);
    p34 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010000001000000000100000000011110",
            TABLE => "111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001001010110110100111111111",
            SHIFT => 2,
            B => -65,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p34_in,
            y(0) => p34_out,
            y(1 to 13 - 1) => dummy34
        );


    p35_in <= x(40) & x(98) & x(198) & x(208) & x(213) & x(256) & x(306) & x(310) & x(338) & x(341) & x(342) & x(343) & x(352) & x(369) & x(370) & x(371) & x(405) & x(415) & x(418) & x(443) & x(446) & x(450) & x(463) & x(471) & x(473) & x(495) & x(497) & x(498) & x(501) & x(522) & x(523) & x(525) & x(552) & x(697);
    y(35) <= not(p35_out);
    p35 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101101001110111010101010111011110",
            TABLE => "0000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101100000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010000001000101011010000100010101110010110011010010000000000000000",
            SHIFT => 2,
            B => 27,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p35_in,
            y(0) => p35_out,
            y(1 to 13 - 1) => dummy35
        );


    p36_in <= x(91) & x(94) & x(118) & x(121) & x(122) & x(134) & x(135) & x(149) & x(171) & x(249) & x(250) & x(276) & x(277) & x(287) & x(304) & x(305) & x(306) & x(329) & x(330) & x(331) & x(342) & x(343) & x(357) & x(358) & x(359) & x(360) & x(362) & x(369) & x(370) & x(371) & x(377) & x(386) & x(387) & x(388) & x(390) & x(391) & x(396) & x(397) & x(416) & x(418) & x(443) & x(473) & x(474) & x(475) & x(501) & x(502) & x(528) & x(529) & x(534) & x(557) & x(584) & x(668) & x(696) & x(697) & x(705) & x(712) & x(713) & x(717) & x(718) & x(720) & x(721) & x(744) & x(745) & x(747) & x(748) & x(749) & x(750);
    y(36) <= not(p36_out);
    p36 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000011000000100011111111101110111001110100000001000000000000000000",
            TABLE => "1111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101101110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 2,
            B => -100,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p36_in,
            y(0) => p36_out,
            y(1 to 14 - 1) => dummy36
        );


    p37_in <= x(66) & x(100) & x(124) & x(125) & x(127) & x(128) & x(136) & x(165) & x(174) & x(179) & x(192) & x(199) & x(220) & x(221) & x(228) & x(248) & x(249) & x(250) & x(256) & x(276) & x(277) & x(278) & x(297) & x(298) & x(299) & x(304) & x(305) & x(306) & x(309) & x(310) & x(311) & x(325) & x(326) & x(333) & x(334) & x(338) & x(339) & x(366) & x(377) & x(405) & x(407) & x(433) & x(473) & x(474) & x(475) & x(557) & x(708) & x(724);
    y(37) <= not(p37_out);
    p37 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011111001101001000100011100011111001110000111110",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p37_in,
            y(0) => p37_out,
            y(1 to 14 - 1) => dummy37
        );


    p38_in <= x(106) & x(133) & x(134) & x(135) & x(136) & x(148) & x(162) & x(163) & x(183) & x(190) & x(191) & x(192) & x(218) & x(220) & x(221) & x(228) & x(248) & x(249) & x(276) & x(277) & x(296) & x(297) & x(298) & x(299) & x(304) & x(305) & x(328) & x(329) & x(330) & x(331) & x(332) & x(358) & x(359) & x(360) & x(361) & x(366) & x(387) & x(388) & x(389) & x(391) & x(396) & x(485) & x(513) & x(717) & x(745);
    y(38) <= not(p38_out);
    p38 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000001001000000100001111001111111111111101111",
            TABLE => "111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => 2,
            B => -19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p38_in,
            y(0) => p38_out,
            y(1 to 13 - 1) => dummy38
        );


    p39_in <= x(44) & x(65) & x(66) & x(67) & x(68) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(191) & x(192) & x(219) & x(247) & x(248) & x(249) & x(276) & x(277) & x(305) & x(328) & x(329) & x(330) & x(331) & x(332) & x(357) & x(358) & x(359) & x(360) & x(361) & x(370) & x(375) & x(376) & x(387) & x(388) & x(389) & x(398) & x(418) & x(514) & x(542) & x(675) & x(707) & x(720) & x(735) & x(736) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(774);
    y(39) <= not(p39_out);
    p39 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000011111111100000000001110001000100000000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 3,
            B => -168,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p39_in,
            y(0) => p39_out,
            y(1 to 14 - 1) => dummy39
        );


    p40_in <= x(65) & x(66) & x(67) & x(68) & x(69) & x(93) & x(198) & x(220) & x(221) & x(247) & x(248) & x(249) & x(250) & x(276) & x(277) & x(289) & x(302) & x(305) & x(306) & x(329) & x(330) & x(331) & x(332) & x(358) & x(359) & x(360) & x(366) & x(369) & x(370) & x(387) & x(424) & x(425) & x(473) & x(501) & x(528) & x(529) & x(600) & x(630);
    y(40) <= not(p40_out);
    p40 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000001001111111011111000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 3,
            B => -86,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p40_in,
            y(0) => p40_out,
            y(1 to 14 - 1) => dummy40
        );


    p41_in <= x(247) & x(248) & x(249) & x(276) & x(277) & x(294) & x(304) & x(305) & x(306) & x(310) & x(329) & x(330) & x(331) & x(333) & x(338) & x(339) & x(357) & x(358) & x(359) & x(360) & x(362) & x(385) & x(386) & x(387) & x(388) & x(486) & x(678) & x(679) & x(705) & x(709) & x(712) & x(717) & x(718) & x(719) & x(739) & x(743) & x(745) & x(746) & x(747);
    y(41) <= not(p41_out);
    p41 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000000011100011110111110000000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 3,
            B => -112,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p41_in,
            y(0) => p41_out,
            y(1 to 14 - 1) => dummy41
        );


    p42_in <= x(106) & x(201) & x(211) & x(228) & x(235) & x(249) & x(256) & x(263) & x(277) & x(283) & x(294) & x(295) & x(296) & x(304) & x(305) & x(306) & x(310) & x(311) & x(321) & x(322) & x(330) & x(333) & x(334) & x(339) & x(357) & x(358) & x(359) & x(360) & x(366) & x(418) & x(474) & x(485) & x(486) & x(487) & x(502) & x(508) & x(514) & x(515) & x(659) & x(695) & x(732) & x(733) & x(769);
    y(42) <= not(p42_out);
    p42 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010000000000000000010001111000111001101110",
            TABLE => "1000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 2,
            B => -70,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p42_in,
            y(0) => p42_out,
            y(1 to 13 - 1) => dummy42
        );


    p43_in <= x(71) & x(106) & x(107) & x(109) & x(165) & x(171) & x(188) & x(189) & x(190) & x(192) & x(194) & x(211) & x(216) & x(217) & x(218) & x(221) & x(243) & x(244) & x(245) & x(246) & x(248) & x(249) & x(266) & x(273) & x(274) & x(276) & x(277) & x(293) & x(294) & x(295) & x(296) & x(303) & x(304) & x(305) & x(306) & x(311) & x(320) & x(321) & x(327) & x(330) & x(331) & x(339) & x(353) & x(354) & x(355) & x(357) & x(358) & x(359) & x(360) & x(366) & x(381) & x(387) & x(390) & x(408) & x(418) & x(435) & x(436) & x(446) & x(451) & x(452) & x(459) & x(463) & x(474) & x(479) & x(480) & x(486) & x(487) & x(502) & x(508) & x(509) & x(510) & x(514) & x(515) & x(516) & x(528) & x(536) & x(537) & x(564) & x(565) & x(566) & x(592) & x(596) & x(620) & x(625) & x(676) & x(704);
    y(43) <= not(p43_out);
    p43 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11100000000100000000000000000000000000111011111110110101100011000110000111000000000000",
            TABLE => "000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 1,
            B => -102,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p43_in,
            y(0) => p43_out,
            y(1 to 13 - 1) => dummy43
        );


    p44_in <= x(35) & x(40) & x(46) & x(49) & x(50) & x(63) & x(64) & x(66) & x(91) & x(108) & x(135) & x(160) & x(186) & x(187) & x(228) & x(257) & x(276) & x(277) & x(301) & x(305) & x(330) & x(331) & x(332) & x(350) & x(359) & x(360) & x(361) & x(378) & x(390) & x(437) & x(446) & x(454) & x(485) & x(571) & x(598) & x(723);
    y(44) <= not(p44_out);
    p44 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111111110011010001000100000111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => 46,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p44_in,
            y(0) => p44_out,
            y(1 to 14 - 1) => dummy44
        );


    p45_in <= x(91) & x(97) & x(98) & x(118) & x(133) & x(134) & x(135) & x(136) & x(160) & x(163) & x(174) & x(187) & x(192) & x(202) & x(221) & x(228) & x(248) & x(249) & x(271) & x(276) & x(277) & x(284) & x(298) & x(299) & x(305) & x(327) & x(328) & x(329) & x(330) & x(331) & x(332) & x(339) & x(351) & x(359) & x(360) & x(361) & x(377) & x(379) & x(387) & x(388) & x(389) & x(390) & x(391) & x(405) & x(406) & x(418) & x(425) & x(473) & x(474) & x(475) & x(502) & x(527) & x(541) & x(555) & x(557) & x(619) & x(688) & x(694) & x(695) & x(705) & x(720) & x(723) & x(732) & x(733);
    y(45) <= not(p45_out);
    p45 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000111111011010110110001000000010001100000110000000000001111111",
            TABLE => "1111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010011000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101101000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 2,
            B => -50,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p45_in,
            y(0) => p45_out,
            y(1 to 14 - 1) => dummy45
        );


    p46_in <= x(66) & x(73) & x(162) & x(163) & x(191) & x(192) & x(220) & x(221) & x(248) & x(249) & x(276) & x(277) & x(304) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(333) & x(346) & x(358) & x(359) & x(360) & x(411) & x(434) & x(438) & x(439) & x(453) & x(454) & x(455) & x(461) & x(466) & x(472) & x(483) & x(484) & x(485) & x(659);
    y(46) <= not(p46_out);
    p46 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000011110011110111110101110",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 2,
            B => -35,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p46_in,
            y(0) => p46_out,
            y(1 to 13 - 1) => dummy46
        );


    p47_in <= x(106) & x(116) & x(304) & x(305) & x(306) & x(313) & x(340) & x(341) & x(342) & x(343) & x(354) & x(368) & x(369) & x(370) & x(377) & x(389) & x(390) & x(391) & x(396) & x(418) & x(446) & x(474) & x(480) & x(485) & x(502) & x(508) & x(509) & x(547) & x(564) & x(767);
    y(47) <= not(p47_out);
    p47 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110001111111110000100001000000",
            TABLE => "010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => -47,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p47_in,
            y(0) => p47_out,
            y(1 to 14 - 1) => dummy47
        );


    p48_in <= x(96) & x(228) & x(248) & x(256) & x(276) & x(277) & x(284) & x(295) & x(304) & x(305) & x(330) & x(331) & x(332) & x(358) & x(359) & x(360) & x(387) & x(388) & x(402) & x(404) & x(405) & x(406) & x(422) & x(431) & x(432) & x(450) & x(507) & x(611) & x(638) & x(639) & x(666) & x(682) & x(694) & x(732);
    y(48) <= not(p48_out);
    p48 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101001000111111110000100110000100",
            TABLE => "0000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101100111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101101000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010011000111000001000100011100001100010010110011010010000000000000000",
            SHIFT => 3,
            B => 20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p48_in,
            y(0) => p48_out,
            y(1 to 14 - 1) => dummy48
        );


    p49_in <= x(35) & x(40) & x(41) & x(46) & x(47) & x(48) & x(50) & x(63) & x(64) & x(66) & x(68) & x(69) & x(70) & x(74) & x(75) & x(78) & x(91) & x(106) & x(107) & x(135) & x(147) & x(173) & x(174) & x(200) & x(201) & x(211) & x(228) & x(229) & x(256) & x(273) & x(274) & x(276) & x(283) & x(299) & x(301) & x(302) & x(305) & x(310) & x(311) & x(338) & x(339) & x(349) & x(359) & x(387) & x(390) & x(396) & x(411) & x(418) & x(423) & x(424) & x(426) & x(446) & x(453) & x(465) & x(466) & x(474) & x(475) & x(491) & x(502) & x(509) & x(531) & x(543) & x(557) & x(558) & x(684) & x(695) & x(723) & x(773) & x(774);
    y(49) <= not(p49_out);
    p49 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000000000000000001111101111101111111110001111111111111111101100011",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 3,
            B => 58,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p49_in,
            y(0) => p49_out,
            y(1 to 15 - 1) => dummy49
        );


    p50_in <= x(171) & x(266) & x(267) & x(268) & x(283) & x(294) & x(295) & x(296) & x(310) & x(311) & x(316) & x(338) & x(339) & x(342) & x(343) & x(349) & x(350) & x(357) & x(358) & x(359) & x(366) & x(370) & x(386) & x(387) & x(389) & x(390) & x(391) & x(418) & x(446) & x(450) & x(473) & x(474) & x(475) & x(501) & x(502) & x(529) & x(557) & x(558) & x(676) & x(690) & x(691) & x(695) & x(705) & x(707) & x(708) & x(709) & x(774);
    y(50) <= not(p50_out);
    p50 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000001001111111011100000000000000011100000",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011000000001000101110001011101111111000000000000000100000001000101111000000100010111000101110111111011101000100000011000000100010111011010011001011010010110011010011001011001101001011010011001011000000001000000000001011100000001000101110000000101111111000101111000000111101000000101111000000100010111100000010111111000010111011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100101111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 2,
            B => -91,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p50_in,
            y(0) => p50_out,
            y(1 to 13 - 1) => dummy50
        );


    p51_in <= x(80) & x(95) & x(96) & x(97) & x(122) & x(126) & x(127) & x(163) & x(164) & x(183) & x(189) & x(190) & x(191) & x(192) & x(194) & x(198) & x(217) & x(218) & x(220) & x(221) & x(222) & x(248) & x(249) & x(276) & x(277) & x(298) & x(304) & x(305) & x(306) & x(326) & x(328) & x(329) & x(330) & x(333) & x(334) & x(338) & x(346) & x(366) & x(370) & x(418) & x(430) & x(458) & x(484) & x(485) & x(507) & x(514) & x(653) & x(720) & x(742) & x(745) & x(746);
    y(51) <= not(p51_out);
    p51 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000011011111011111111101110000110101000001010000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 2,
            B => 38,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p51_in,
            y(0) => p51_out,
            y(1 to 13 - 1) => dummy51
        );


    p52_in <= x(67) & x(89) & x(90) & x(91) & x(92) & x(93) & x(94) & x(193) & x(250) & x(274) & x(303) & x(307) & x(330) & x(331) & x(332) & x(358) & x(359) & x(360) & x(361) & x(387) & x(389) & x(396) & x(479) & x(480) & x(507) & x(537) & x(564) & x(565) & x(567) & x(593) & x(594) & x(619) & x(622) & x(638) & x(647) & x(666) & x(688);
    y(52) <= not(p52_out);
    p52 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000000000000000001000000000001010",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => -170,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p52_in,
            y(0) => p52_out,
            y(1 to 14 - 1) => dummy52
        );


    p53_in <= x(106) & x(134) & x(135) & x(147) & x(163) & x(174) & x(176) & x(203) & x(204) & x(205) & x(206) & x(230) & x(231) & x(234) & x(235) & x(257) & x(258) & x(269) & x(272) & x(285) & x(286) & x(295) & x(300) & x(301) & x(302) & x(313) & x(327) & x(330) & x(332) & x(360) & x(361) & x(362) & x(366) & x(389) & x(390) & x(391) & x(418) & x(446) & x(451) & x(474) & x(475) & x(479) & x(531) & x(555) & x(707);
    y(53) <= not(p53_out);
    p53 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111010000000000000000100000000000000000000000",
            TABLE => "000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 2,
            B => -116,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p53_in,
            y(0) => p53_out,
            y(1 to 13 - 1) => dummy53
        );


    p54_in <= x(248) & x(267) & x(276) & x(277) & x(278) & x(305) & x(306) & x(329) & x(330) & x(331) & x(333) & x(334) & x(358) & x(359) & x(360) & x(379) & x(380) & x(387) & x(388) & x(397) & x(398) & x(399) & x(415) & x(416) & x(424) & x(425) & x(426) & x(443) & x(453) & x(454) & x(553) & x(558) & x(564) & x(619) & x(649) & x(691) & x(697) & x(707) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(748) & x(750);
    y(54) <= not(p54_out);
    p54 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10111110001100011000000000000000000101111111111",
            TABLE => "00000001000101110000000000000001000101110111111100000001000101111000000100010111111010001000000100010111011111101000000100010111011010011001011010010110011010011001011001101001011010011001011001110001000100000001000000000000111101110111000101110001000100000111000100011000000110001000111011100111011100010111000100011000011010011001011010010110011010011001011001101001011010011001011010111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111101110101001101010001000000110101000100000001000000000000001011110111010100110101000100001011010100010000100100001000101011011010011001011010010110011010011001011001101001011010011001011000000001000101110001011101111111000000000000000100000001000101111000000100010111000101110111111011101000100000011000000100010111011010011001011010010110011010011001011001101001011010011001011000000001000101110001011101111111100000010001011100010111011111100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 2,
            B => -26,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p54_in,
            y(0) => p54_out,
            y(1 to 13 - 1) => dummy54
        );


    p55_in <= x(128) & x(156) & x(157) & x(158) & x(165) & x(192) & x(221) & x(249) & x(250) & x(274) & x(277) & x(305) & x(306) & x(331) & x(333) & x(334) & x(359) & x(360) & x(387) & x(388) & x(390) & x(418) & x(450) & x(451) & x(474) & x(480) & x(508) & x(509) & x(510) & x(520) & x(536) & x(537) & x(539) & x(540) & x(541) & x(547) & x(554) & x(564) & x(565) & x(566) & x(567) & x(568) & x(582) & x(583) & x(584) & x(592) & x(593) & x(594) & x(595) & x(609) & x(610) & x(611) & x(620) & x(638) & x(664) & x(665) & x(666);
    y(55) <= not(p55_out);
    p55 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000000000010011110010000000000000000000000000000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 2,
            B => -126,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p55_in,
            y(0) => p55_out,
            y(1 to 13 - 1) => dummy55
        );


    p56_in <= x(66) & x(220) & x(247) & x(248) & x(275) & x(276) & x(277) & x(306) & x(317) & x(453) & x(480) & x(501) & x(502) & x(507) & x(529) & x(535) & x(564) & x(660) & x(705) & x(733);
    y(56) <= not(p56_out);
    p56 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111100000000100",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p56_in,
            y(0) => p56_out,
            y(1 to 14 - 1) => dummy56
        );


    p57_in <= x(64) & x(66) & x(70) & x(71) & x(108) & x(136) & x(145) & x(165) & x(171) & x(192) & x(221) & x(241) & x(248) & x(249) & x(256) & x(272) & x(273) & x(274) & x(276) & x(277) & x(283) & x(301) & x(302) & x(305) & x(306) & x(310) & x(311) & x(333) & x(334) & x(339) & x(358) & x(359) & x(360) & x(366) & x(378) & x(387) & x(403) & x(404) & x(406) & x(422) & x(431) & x(432) & x(445) & x(459) & x(473) & x(486) & x(574) & x(602) & x(603) & x(675) & x(676) & x(677) & x(679) & x(697) & x(704) & x(705) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(713);
    y(57) <= not(p57_out);
    p57 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111100000000000000000000000001110111110111111111000010000000000",
            TABLE => "0000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011101010001000000010000000000000011111101110101001101010001000000110101000100001001000010001010111011110111010100110101000100001010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 2,
            B => -104,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p57_in,
            y(0) => p57_out,
            y(1 to 14 - 1) => dummy57
        );


    p58_in <= x(122) & x(176) & x(178) & x(242) & x(269) & x(350) & x(351) & x(354) & x(377) & x(381) & x(433) & x(435) & x(490) & x(501) & x(502) & x(529) & x(557) & x(742) & x(746);
    y(58) <= not(p58_out);
    p58 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000011111111000000",
            TABLE => "1111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 3,
            B => -40,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p58_in,
            y(0) => p58_out,
            y(1 to 13 - 1) => dummy58
        );


    p59_in <= x(136) & x(320) & x(321) & x(333) & x(340) & x(341) & x(342) & x(343) & x(369) & x(401) & x(402) & x(422) & x(427) & x(428) & x(429) & x(454) & x(473) & x(501) & x(528) & x(529) & x(583) & x(611) & x(697) & x(705) & x(707) & x(709) & x(713) & x(714) & x(715) & x(716) & x(717) & x(719) & x(720) & x(721) & x(722) & x(744) & x(746) & x(747) & x(748) & x(750);
    y(59) <= not(p59_out);
    p59 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111111110010000000000011111111111111111",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 3,
            B => 80,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p59_in,
            y(0) => p59_out,
            y(1 to 14 - 1) => dummy59
        );


    p60_in <= x(44) & x(65) & x(66) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(91) & x(93) & x(94) & x(97) & x(99) & x(100) & x(233) & x(234) & x(277) & x(330) & x(331) & x(338) & x(342) & x(343) & x(348) & x(349) & x(358) & x(359) & x(360) & x(366) & x(369) & x(370) & x(371) & x(387) & x(397) & x(417) & x(418) & x(446) & x(473) & x(474) & x(492) & x(493) & x(501) & x(517) & x(528) & x(529) & x(541) & x(739) & x(742) & x(743) & x(744) & x(745) & x(750);
    y(60) <= not(p60_out);
    p60 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111111111111110010010000000100000111110011111111111",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010011110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101101111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101101111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 2,
            B => 114,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p60_in,
            y(0) => p60_out,
            y(1 to 13 - 1) => dummy60
        );


    p61_in <= x(35) & x(46) & x(62) & x(63) & x(66) & x(68) & x(69) & x(70) & x(73) & x(74) & x(75) & x(76) & x(78) & x(79) & x(91) & x(93) & x(94) & x(95) & x(96) & x(97) & x(101) & x(102) & x(103) & x(104) & x(106) & x(107) & x(108) & x(146) & x(171) & x(199) & x(206) & x(228) & x(248) & x(255) & x(256) & x(275) & x(276) & x(277) & x(305) & x(310) & x(311) & x(338) & x(339) & x(366) & x(376) & x(403) & x(404) & x(445) & x(450) & x(535) & x(563) & x(649) & x(676) & x(677) & x(678) & x(679) & x(680) & x(691) & x(704) & x(705) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(714) & x(715) & x(736) & x(750);
    y(61) <= not(p61_out);
    p61 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111111111111111111111111111011000011111000111111111101111111111111",
            TABLE => "00000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000010000000000010101100000010001010110000001010111111001010110100001011010100001010110100001000101011010000101011110100101011100101100110100101101001100101100110100110010110100101100110100101111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011001000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000100000001000001110001000100000111000101110001111101111000111000011000000110000111000100011000011100010111000111100111011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000001000101110001011101111111100000010001011100010111011111100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 3,
            B => 415,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p61_in,
            y(0) => p61_out,
            y(1 to 15 - 1) => dummy61
        );


    p62_in <= x(35) & x(41) & x(44) & x(64) & x(124) & x(133) & x(151) & x(152) & x(305) & x(331) & x(332) & x(338) & x(339) & x(357) & x(358) & x(359) & x(360) & x(366) & x(385) & x(386) & x(387) & x(388) & x(391) & x(414) & x(415) & x(416) & x(418) & x(446) & x(474) & x(475) & x(529) & x(531) & x(584) & x(696) & x(750);
    y(62) <= not(p62_out);
    p62 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11010100011001111011110111000000000",
            TABLE => "00000100000000000100110100000100010011010000010011011111010011010010010010110010010011010010010001001101001001001101101101001101100101100110100101101001100101100110100110010110100101100110100110111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100100000010001010110010101110111111000000000000001000000010001010110100001000101011001010111011110111010100010000100100001000101011100101100110100101101001100101100110100110010110100101100110100100000000000001000000010001001101000001000100110101001101110111111011001000100100001001000100110100100100010011010100110111011011011010011001011010010110011010011001011001101001011010011001011010000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p62_in,
            y(0) => p62_out,
            y(1 to 14 - 1) => dummy62
        );


    p63_in <= x(117) & x(248) & x(249) & x(276) & x(277) & x(303) & x(304) & x(305) & x(306) & x(322) & x(333) & x(334) & x(359) & x(360) & x(387) & x(388) & x(455) & x(501) & x(707) & x(718) & x(719) & x(720) & x(742) & x(745) & x(746);
    y(63) <= not(p63_out);
    p63 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000000000001111110000000",
            TABLE => "1110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -159,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p63_in,
            y(0) => p63_out,
            y(1 to 14 - 1) => dummy63
        );


    p64_in <= x(35) & x(64) & x(78) & x(106) & x(107) & x(192) & x(217) & x(218) & x(220) & x(221) & x(243) & x(244) & x(245) & x(246) & x(248) & x(249) & x(273) & x(274) & x(276) & x(277) & x(305) & x(306) & x(322) & x(330) & x(331) & x(334) & x(341) & x(347) & x(350) & x(357) & x(358) & x(359) & x(360) & x(369) & x(375) & x(386) & x(387) & x(390) & x(415) & x(418) & x(446) & x(465) & x(473) & x(474) & x(501) & x(502) & x(528) & x(635) & x(637) & x(719) & x(720) & x(721) & x(742) & x(746);
    y(64) <= not(p64_out);
    p64 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000001111111111111111100010100000010010111111111100000",
            TABLE => "111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 2,
            B => 25,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p64_in,
            y(0) => p64_out,
            y(1 to 13 - 1) => dummy64
        );


    p65_in <= x(35) & x(46) & x(62) & x(63) & x(64) & x(66) & x(68) & x(69) & x(70) & x(78) & x(90) & x(91) & x(103) & x(104) & x(107) & x(108) & x(249) & x(250) & x(277) & x(278) & x(305) & x(306) & x(338) & x(396) & x(424) & x(450) & x(507) & x(521) & x(549) & x(557) & x(576) & x(578) & x(591) & x(605) & x(634) & x(647) & x(662) & x(676) & x(683) & x(684) & x(685) & x(686) & x(687) & x(688);
    y(65) <= not(p65_out);
    p65 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111111111111111110001111011111111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 3,
            B => 186,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p65_in,
            y(0) => p65_out,
            y(1 to 14 - 1) => dummy65
        );


    p66_in <= x(64) & x(72) & x(91) & x(92) & x(93) & x(95) & x(108) & x(315) & x(341) & x(342) & x(355) & x(360) & x(369) & x(382) & x(387) & x(388) & x(389) & x(416) & x(417) & x(473) & x(501) & x(527) & x(528) & x(529) & x(619) & x(720);
    y(66) <= not(p66_out);
    p66 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01000001111011000000000001",
            TABLE => "111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 3,
            B => -139,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p66_in,
            y(0) => p66_out,
            y(1 to 13 - 1) => dummy66
        );


    p67_in <= x(177) & x(192) & x(220) & x(221) & x(237) & x(238) & x(248) & x(249) & x(266) & x(267) & x(268) & x(275) & x(276) & x(277) & x(294) & x(295) & x(296) & x(305) & x(309) & x(323) & x(338) & x(343) & x(366) & x(370) & x(371) & x(398) & x(399) & x(418) & x(473) & x(474) & x(501) & x(502) & x(664) & x(665) & x(718) & x(739) & x(742) & x(744) & x(747);
    y(67) <= not(p67_out);
    p67 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000011001110001110111010000111110011111",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 2,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p67_in,
            y(0) => p67_out,
            y(1 to 13 - 1) => dummy67
        );


    p68_in <= x(95) & x(98) & x(117) & x(118) & x(121) & x(122) & x(124) & x(125) & x(126) & x(127) & x(128) & x(133) & x(135) & x(147) & x(148) & x(149) & x(152) & x(163) & x(191) & x(192) & x(220) & x(221) & x(248) & x(249) & x(266) & x(267) & x(276) & x(277) & x(302) & x(304) & x(305) & x(306) & x(318) & x(328) & x(329) & x(330) & x(331) & x(332) & x(346) & x(357) & x(358) & x(359) & x(360) & x(387) & x(389) & x(453) & x(474) & x(475) & x(502) & x(613) & x(619) & x(736) & x(738) & x(746);
    y(68) <= not(p68_out);
    p68 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111110011110000000110010000111110111111111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 2,
            B => 68,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p68_in,
            y(0) => p68_out,
            y(1 to 13 - 1) => dummy68
        );


    p69_in <= x(182) & x(210) & x(211) & x(232) & x(233) & x(234) & x(238) & x(260) & x(269) & x(270) & x(276) & x(310) & x(329) & x(338) & x(339) & x(350) & x(357) & x(366) & x(378) & x(406) & x(407) & x(440) & x(467) & x(469) & x(494) & x(501) & x(518) & x(528) & x(695) & x(704) & x(719) & x(720) & x(738);
    y(69) <= not(p69_out);
    p69 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111000100000100110111000001010111",
            TABLE => "000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 2,
            B => -37,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p69_in,
            y(0) => p69_out,
            y(1 to 13 - 1) => dummy69
        );


    p70_in <= x(97) & x(100) & x(127) & x(135) & x(136) & x(155) & x(156) & x(163) & x(164) & x(192) & x(194) & x(213) & x(221) & x(222) & x(248) & x(249) & x(276) & x(277) & x(305) & x(328) & x(329) & x(330) & x(331) & x(332) & x(338) & x(356) & x(357) & x(358) & x(359) & x(360) & x(361) & x(368) & x(370) & x(387) & x(388) & x(389) & x(390) & x(391) & x(396) & x(418) & x(474) & x(484) & x(485) & x(512) & x(513) & x(535) & x(547) & x(575) & x(675) & x(676) & x(705) & x(706) & x(710) & x(711) & x(712) & x(713) & x(723) & x(745) & x(746);
    y(70) <= not(p70_out);
    p70 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00011001111111111110000000000001100000100000010011111111100",
            TABLE => "10111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100100000001000101110001011101111111000000000000000100000001000101111000000100010111000101110111111011101000100000011000000100010111011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100111101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100110000000111010001110100011111110000000001000000010000000111010001000000111101000111010000111111000010111100000011000000111101000100101100110100101101001100101100110100110010110100101100110100111101000111111101000000011101000100000001110100000000000100000001110100001111110100000011110100010000001111010000001011110000001011010011001011010010110011010011001011001101001011010011001011011101111100011101000111000001000100011100000100000001000000000001110011110001110100011100001100010001110000110000001100001110001011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100001000100011101000111011101111000110001000111010001110111001110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 2,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p70_in,
            y(0) => p70_out,
            y(1 to 14 - 1) => dummy70
        );


    p71_in <= x(35) & x(41) & x(78) & x(133) & x(135) & x(202) & x(230) & x(256) & x(257) & x(270) & x(273) & x(274) & x(285) & x(311) & x(321) & x(322) & x(349) & x(350) & x(351) & x(358) & x(369) & x(389) & x(390) & x(446) & x(473) & x(502) & x(507) & x(509) & x(535) & x(637) & x(664) & x(695) & x(720) & x(746) & x(769);
    y(71) <= not(p71_out);
    p71 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000111111111000000011111111110001",
            TABLE => "11111101110101001101010001000000110101000100000001000000000000001011110111010100110101000100001011010100010000100100001000101011011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100110000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100101111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100111010100010000001111110111010100110101000100001010111101110101001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => 51,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p71_in,
            y(0) => p71_out,
            y(1 to 14 - 1) => dummy71
        );


    p72_in <= x(39) & x(40) & x(41) & x(46) & x(159) & x(160) & x(186) & x(187) & x(188) & x(192) & x(198) & x(200) & x(214) & x(228) & x(248) & x(249) & x(257) & x(275) & x(276) & x(277) & x(303) & x(304) & x(305) & x(306) & x(324) & x(328) & x(330) & x(333) & x(334) & x(338) & x(366) & x(381) & x(437) & x(464) & x(465) & x(491) & x(518) & x(528) & x(570) & x(655) & x(681) & x(724) & x(741) & x(742) & x(774);
    y(72) <= not(p72_out);
    p72 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111100101101111111000110000000011111000",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 2,
            B => 56,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p72_in,
            y(0) => p72_out,
            y(1 to 13 - 1) => dummy72
        );


    p73_in <= x(215) & x(216) & x(242) & x(243) & x(244) & x(249) & x(266) & x(277) & x(294) & x(295) & x(305) & x(309) & x(310) & x(312) & x(314) & x(322) & x(333) & x(338) & x(339) & x(358) & x(359) & x(360) & x(366) & x(387) & x(388) & x(403) & x(427) & x(429) & x(456) & x(458) & x(459) & x(484) & x(486) & x(501) & x(512) & x(623) & x(625) & x(651) & x(665) & x(666) & x(677) & x(679) & x(707) & x(708) & x(709) & x(711) & x(712) & x(713) & x(714) & x(715) & x(737) & x(744) & x(750);
    y(73) <= not(p73_out);
    p73 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000000001110111111111111000110000000000000",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000100000001000101011000000100010101100101011101111111101010001000010010000100010101101000010001010110010101110111101011010011001011010010110011010011001011001101001011010011001011010001110111011110000100010001110000010001000111000000000000010001000111011100111000110001000111000011000100011100111000100011000100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 2,
            B => -72,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p73_in,
            y(0) => p73_out,
            y(1 to 13 - 1) => dummy73
        );


    p74_in <= x(248) & x(249) & x(276) & x(277) & x(305) & x(306) & x(330) & x(357) & x(358) & x(359) & x(360) & x(388) & x(424) & x(425) & x(428) & x(453) & x(659) & x(704) & x(705) & x(750);
    y(74) <= not(p74_out);
    p74 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111100000000001111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 3,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p74_in,
            y(0) => p74_out,
            y(1 to 13 - 1) => dummy74
        );


    p75_in <= x(65) & x(66) & x(93) & x(94) & x(118) & x(124) & x(190) & x(192) & x(198) & x(219) & x(220) & x(221) & x(247) & x(248) & x(249) & x(275) & x(276) & x(277) & x(294) & x(303) & x(304) & x(305) & x(306) & x(347) & x(371) & x(372) & x(373) & x(374) & x(375) & x(400) & x(413) & x(414) & x(415) & x(416) & x(434) & x(440) & x(442) & x(443) & x(450) & x(461) & x(468) & x(475) & x(485) & x(486) & x(488) & x(513) & x(583) & x(613) & x(654) & x(666) & x(675) & x(717) & x(737) & x(739) & x(740) & x(742) & x(744) & x(745) & x(746);
    y(75) <= not(p75_out);
    p75 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000011011111111101111111111111110111101000000010100000000",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100000001000000000001011100000001000101110000000101111111000101111000000111101000000101111000000100010111100000010111111000010111011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000001000101110001011101111111000000000000000100000001000101111000000100010111000101110111111011101000100000011000000100010111011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000001000000010001001101000001000100110101001101110111111011001000100100001001000100110100100100010011010100110111011011011010011001011010010110011010011001011001101001011010011001011000000000001000000010000010110010001000001011001010110010111110110100110100100100001001001011001000100100101100101011001011011011100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100110000000111010000000000010000000111010001111111010000000111010001000000111101000000101111000000111101000011111101000000111101000100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 2,
            B => 24,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p75_in,
            y(0) => p75_out,
            y(1 to 14 - 1) => dummy75
        );


    p76_in <= x(44) & x(118) & x(135) & x(163) & x(191) & x(192) & x(200) & x(219) & x(220) & x(221) & x(228) & x(247) & x(248) & x(249) & x(275) & x(276) & x(277) & x(304) & x(305) & x(306) & x(318) & x(327) & x(328) & x(329) & x(330) & x(342) & x(343) & x(344) & x(346) & x(347) & x(348) & x(349) & x(350) & x(355) & x(360) & x(361) & x(369) & x(370) & x(371) & x(373) & x(374) & x(379) & x(389) & x(390) & x(391) & x(417) & x(418) & x(443) & x(446) & x(453) & x(454) & x(473) & x(474) & x(475) & x(480) & x(502);
    y(76) <= not(p76_out);
    p76 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00111101110111111111100001111111100011111100000100000000",
            TABLE => "000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 2,
            B => 18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p76_in,
            y(0) => p76_out,
            y(1 to 13 - 1) => dummy76
        );


    p77_in <= x(35) & x(63) & x(91) & x(108) & x(161) & x(162) & x(190) & x(191) & x(209) & x(210) & x(211) & x(212) & x(330) & x(339) & x(355) & x(356) & x(367) & x(379) & x(485) & x(486) & x(528) & x(543) & x(544) & x(603) & x(605) & x(632) & x(659) & x(695) & x(719) & x(720);
    y(77) <= not(p77_out);
    p77 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111110000010010001111111000",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => 52,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p77_in,
            y(0) => p77_out,
            y(1 to 14 - 1) => dummy77
        );


    p78_in <= x(106) & x(123) & x(210) & x(211) & x(212) & x(220) & x(231) & x(248) & x(249) & x(276) & x(277) & x(305) & x(310) & x(312) & x(331) & x(338) & x(339) & x(340) & x(349) & x(358) & x(359) & x(360) & x(366) & x(376) & x(387) & x(416) & x(425) & x(438) & x(453) & x(538) & x(553) & x(581) & x(707);
    y(78) <= not(p78_out);
    p78 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100001111111110111000010000100001",
            TABLE => "110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110110101001001011011111111",
            SHIFT => 3,
            B => 15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p78_in,
            y(0) => p78_out,
            y(1 to 14 - 1) => dummy78
        );


    p79_in <= x(48) & x(50) & x(91) & x(182) & x(221) & x(248) & x(293) & x(294) & x(295) & x(296) & x(305) & x(310) & x(321) & x(322) & x(338) & x(339) & x(366) & x(375) & x(424) & x(501) & x(553) & x(606) & x(611) & x(637) & x(638) & x(639) & x(665) & x(666) & x(667) & x(694) & x(695) & x(707) & x(708) & x(709) & x(710) & x(711) & x(715) & x(744) & x(745) & x(747) & x(750);
    y(79) <= not(p79_out);
    p79 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00011100001000000111111111111110000000000",
            TABLE => "01111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011011111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011011111101110101001101010001000000110101000100000001000000000000001011110111010100110101000100001011010100010000100100001000101011011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100111101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p79_in,
            y(0) => p79_out,
            y(1 to 14 - 1) => dummy79
        );


    p80_in <= x(44) & x(65) & x(80) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(108) & x(118) & x(119) & x(121) & x(148) & x(163) & x(192) & x(248) & x(249) & x(276) & x(277) & x(305) & x(318) & x(322) & x(323) & x(338) & x(349) & x(350) & x(351) & x(366) & x(369) & x(370) & x(377) & x(378) & x(379) & x(389) & x(391) & x(406) & x(417) & x(418) & x(454) & x(465) & x(473) & x(474) & x(475) & x(482) & x(492) & x(493) & x(501) & x(520) & x(521) & x(522) & x(528) & x(529) & x(549) & x(661) & x(743) & x(770);
    y(80) <= not(p80_out);
    p80 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000000000001111111111011101111100100000000000000000100",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100011101001011011111111",
            SHIFT => 2,
            B => -61,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p80_in,
            y(0) => p80_out,
            y(1 to 13 - 1) => dummy80
        );


    p81_in <= x(95) & x(97) & x(108) & x(192) & x(220) & x(221) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(278) & x(304) & x(305) & x(306) & x(320) & x(321) & x(322) & x(328) & x(329) & x(330) & x(333) & x(334) & x(341) & x(342) & x(343) & x(344) & x(348) & x(349) & x(350) & x(370) & x(371) & x(418) & x(446) & x(473) & x(474) & x(501) & x(502) & x(528) & x(529) & x(557) & x(613) & x(697);
    y(81) <= not(p81_out);
    p81 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000111111111111111110001111111111100000000000",
            TABLE => "011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 3,
            B => 33,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p81_in,
            y(0) => p81_out,
            y(1 to 14 - 1) => dummy81
        );


    p82_in <= x(65) & x(67) & x(93) & x(94) & x(96) & x(97) & x(229) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(305) & x(306) & x(333) & x(334) & x(358) & x(359) & x(360) & x(362) & x(369) & x(370) & x(380) & x(387) & x(388) & x(390) & x(396) & x(397) & x(398) & x(399) & x(418) & x(424) & x(425) & x(433) & x(451) & x(473) & x(474) & x(479) & x(501) & x(529) & x(713) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(744) & x(745) & x(747) & x(748) & x(749) & x(750);
    y(82) <= not(p82_out);
    p82 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000001000000000011101101101111011000000000000000000000",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010010000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100000100010001110000000000000100010001110111011110000100010001110000110001000111001110001000110001000111011100111000110001000111001101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => -220,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p82_in,
            y(0) => p82_out,
            y(1 to 14 - 1) => dummy82
        );


    p83_in <= x(145) & x(207) & x(212) & x(247) & x(248) & x(249) & x(250) & x(276) & x(277) & x(304) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(333) & x(357) & x(358) & x(359) & x(360) & x(366) & x(387) & x(388) & x(390) & x(391) & x(408) & x(418) & x(436) & x(437) & x(446) & x(454) & x(455) & x(473) & x(474) & x(483) & x(500) & x(501) & x(502) & x(528) & x(529) & x(556) & x(557) & x(584) & x(656) & x(747) & x(748) & x(750);
    y(83) <= not(p83_out);
    p83 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011111111111000010000100110100100110111111111111",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => 96,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p83_in,
            y(0) => p83_out,
            y(1 to 14 - 1) => dummy83
        );


    p84_in <= x(136) & x(145) & x(164) & x(171) & x(172) & x(194) & x(221) & x(222) & x(228) & x(305) & x(311) & x(368) & x(369) & x(379) & x(403) & x(407) & x(422) & x(430) & x(431) & x(473) & x(474) & x(535) & x(575) & x(675) & x(676) & x(677) & x(678) & x(679) & x(704) & x(705) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(736);
    y(84) <= not(p84_out);
    p84 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000000000111011110100000000000000",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => -205,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p84_in,
            y(0) => p84_out,
            y(1 to 14 - 1) => dummy84
        );


    p85_in <= x(72) & x(136) & x(178) & x(206) & x(230) & x(247) & x(294) & x(295) & x(305) & x(321) & x(322) & x(323) & x(333) & x(334) & x(340) & x(341) & x(342) & x(343) & x(350) & x(359) & x(360) & x(368) & x(369) & x(387) & x(388) & x(389) & x(403) & x(446) & x(455) & x(458) & x(473) & x(486) & x(501) & x(511) & x(514) & x(516) & x(528) & x(611) & x(653) & x(654) & x(655) & x(658) & x(675) & x(677) & x(679) & x(683) & x(707) & x(708) & x(709) & x(719) & x(745) & x(746);
    y(85) <= not(p85_out);
    p85 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111101111111111111001100000000000000011111111111111",
            TABLE => "0000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 2,
            B => 45,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p85_in,
            y(0) => p85_out,
            y(1 to 13 - 1) => dummy85
        );


    p86_in <= x(185) & x(192) & x(199) & x(219) & x(220) & x(221) & x(228) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(320) & x(328) & x(329) & x(330) & x(333) & x(354) & x(357) & x(358) & x(359) & x(360) & x(388) & x(390) & x(418) & x(434) & x(435) & x(446) & x(487) & x(489) & x(509) & x(510) & x(515) & x(528) & x(611) & x(695);
    y(86) <= not(p86_out);
    p86 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010001000000000000011101111110011011001001",
            TABLE => "1000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010010101110111111000000100010101100000010001010110000000000000010001010111011110101000010001010110100001000101011110101000100001001101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010100110111011111000001000100110100000100010011010000000000000100010011011101101100100100010011010010010001001101101100100010010001101001100101101001011001101001100101100110100101101001100101101000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => -96,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p86_in,
            y(0) => p86_out,
            y(1 to 14 - 1) => dummy86
        );


    p87_in <= x(186) & x(188) & x(214) & x(239) & x(240) & x(244) & x(250) & x(276) & x(277) & x(303) & x(304) & x(305) & x(306) & x(333) & x(334) & x(357) & x(358) & x(359) & x(360) & x(362) & x(367) & x(384) & x(390) & x(391) & x(396) & x(412) & x(418) & x(426) & x(479) & x(480) & x(485) & x(486) & x(508) & x(516) & x(535) & x(537) & x(564) & x(565) & x(592) & x(593) & x(625) & x(635) & x(654) & x(662) & x(676) & x(688) & x(689) & x(696) & x(724) & x(748);
    y(87) <= not(p87_out);
    p87 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111111111100001101100101100101111111111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 2,
            B => 115,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p87_in,
            y(0) => p87_out,
            y(1 to 13 - 1) => dummy87
        );


    p88_in <= x(64) & x(66) & x(78) & x(106) & x(135) & x(144) & x(147) & x(173) & x(174) & x(175) & x(183) & x(185) & x(200) & x(201) & x(202) & x(210) & x(211) & x(212) & x(229) & x(257) & x(276) & x(311) & x(316) & x(342) & x(359) & x(369) & x(379) & x(389) & x(390) & x(407) & x(418) & x(424) & x(446) & x(452) & x(474) & x(475) & x(480) & x(502) & x(557) & x(558) & x(619) & x(649) & x(695) & x(697) & x(718) & x(719) & x(720) & x(721) & x(723) & x(773);
    y(88) <= not(p88_out);
    p88 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111000001100011100101111100100000000000010111110",
            TABLE => "000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 3,
            B => -85,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p88_in,
            y(0) => p88_out,
            y(1 to 14 - 1) => dummy88
        );


    p89_in <= x(100) & x(192) & x(221) & x(238) & x(248) & x(249) & x(266) & x(267) & x(276) & x(277) & x(294) & x(296) & x(305) & x(338) & x(347) & x(366) & x(375) & x(376) & x(418) & x(474) & x(544) & x(545) & x(546) & x(573) & x(574) & x(633) & x(634) & x(653) & x(655) & x(656) & x(657) & x(662) & x(663) & x(681) & x(683) & x(742) & x(744) & x(745) & x(747);
    y(89) <= not(p89_out);
    p89 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100100110011010100111111100000000001111",
            TABLE => "100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => 2,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p89_in,
            y(0) => p89_out,
            y(1 to 13 - 1) => dummy89
        );


    p90_in <= x(44) & x(134) & x(135) & x(165) & x(180) & x(181) & x(236) & x(238) & x(245) & x(250) & x(264) & x(266) & x(274) & x(286) & x(301) & x(333) & x(362) & x(369) & x(370) & x(387) & x(390) & x(391) & x(396) & x(397) & x(398) & x(399) & x(400) & x(401) & x(416) & x(418) & x(429) & x(430) & x(451) & x(474) & x(475) & x(531) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(713) & x(714) & x(715) & x(717) & x(736) & x(737) & x(738) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(750) & x(764);
    y(90) <= not(p90_out);
    p90 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110000000000000011100111111101100000000000000000000000000",
            TABLE => "1000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010010000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 2,
            B => -101,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p90_in,
            y(0) => p90_out,
            y(1 to 14 - 1) => dummy90
        );


    p91_in <= x(65) & x(91) & x(109) & x(137) & x(192) & x(221) & x(248) & x(249) & x(276) & x(277) & x(304) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(332) & x(341) & x(357) & x(358) & x(359) & x(360) & x(361) & x(384) & x(387) & x(388) & x(391) & x(407) & x(418) & x(434) & x(435) & x(473) & x(474) & x(490) & x(494) & x(501) & x(502) & x(508) & x(521) & x(522) & x(523) & x(528) & x(529) & x(557) & x(568) & x(579) & x(584) & x(592) & x(606) & x(611) & x(626) & x(668) & x(696) & x(705) & x(739) & x(742) & x(743) & x(745) & x(766);
    y(91) <= not(p91_out);
    p91 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000000000011111111111111010110010000000000000000000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 2,
            B => -126,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p91_in,
            y(0) => p91_out,
            y(1 to 14 - 1) => dummy91
        );


    p92_in <= x(66) & x(192) & x(221) & x(249) & x(276) & x(277) & x(305) & x(330) & x(331) & x(338) & x(348) & x(349) & x(350) & x(358) & x(360) & x(366) & x(377) & x(389) & x(390) & x(391) & x(418) & x(446) & x(474) & x(501) & x(502) & x(507) & x(514) & x(528) & x(529) & x(675) & x(709) & x(710) & x(720) & x(723);
    y(92) <= not(p92_out);
    p92 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000111000111011111111011100000",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010011110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 3,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p92_in,
            y(0) => p92_out,
            y(1 to 14 - 1) => dummy92
        );


    p93_in <= x(44) & x(165) & x(192) & x(220) & x(221) & x(246) & x(247) & x(248) & x(249) & x(250) & x(273) & x(274) & x(275) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(307) & x(333) & x(334) & x(378) & x(389) & x(390) & x(396) & x(418) & x(443) & x(444) & x(446) & x(451) & x(471) & x(479) & x(486) & x(489) & x(500) & x(526) & x(537) & x(628) & x(655) & x(656) & x(683) & x(724) & x(738);
    y(93) <= not(p93_out);
    p93 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111111111111111110110111111100111111110",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001001010110110100111111111",
            SHIFT => 2,
            B => 163,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p93_in,
            y(0) => p93_out,
            y(1 to 13 - 1) => dummy93
        );


    p94_in <= x(44) & x(91) & x(92) & x(94) & x(96) & x(266) & x(277) & x(294) & x(305) & x(306) & x(310) & x(316) & x(330) & x(333) & x(342) & x(343) & x(357) & x(358) & x(359) & x(360) & x(369) & x(370) & x(371) & x(387) & x(396) & x(397) & x(398) & x(418) & x(426) & x(446) & x(450) & x(473) & x(474) & x(486) & x(501) & x(502) & x(529) & x(676) & x(684) & x(685) & x(718) & x(722) & x(724) & x(750);
    y(94) <= not(p94_out);
    p94 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000110111111111111101000010000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 2,
            B => -45,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p94_in,
            y(0) => p94_out,
            y(1 to 13 - 1) => dummy94
        );


    p95_in <= x(145) & x(171) & x(249) & x(261) & x(262) & x(288) & x(289) & x(315) & x(317) & x(343) & x(344) & x(359) & x(387) & x(388) & x(397) & x(415) & x(416) & x(507) & x(516) & x(528) & x(656) & x(657) & x(742);
    y(95) <= not(p95_out);
    p95 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11100000000000000100111",
            TABLE => "00000000100000001000000011101000100000001110100011101000111111100001011110000001100000011110100010000001111010001110100001111110011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111101110101001101010001000000110101000100000001000000000000001011110111010100110101000100001011010100010000100100001000101011011010011001011010010110011010011001011001101001011010011001011001111111000101110001011100000001011111100001011100010111100000010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 2,
            B => -38,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p95_in,
            y(0) => p95_out,
            y(1 to 12 - 1) => dummy95
        );


    p96_in <= x(107) & x(109) & x(122) & x(124) & x(149) & x(150) & x(151) & x(165) & x(194) & x(210) & x(243) & x(249) & x(277) & x(293) & x(305) & x(321) & x(322) & x(345) & x(348) & x(349) & x(350) & x(359) & x(360) & x(369) & x(387) & x(388) & x(390) & x(391) & x(418) & x(446) & x(473) & x(474) & x(480) & x(481) & x(499) & x(501) & x(502) & x(508) & x(509) & x(510) & x(528) & x(536) & x(537) & x(538) & x(539) & x(550) & x(552) & x(553) & x(554) & x(557) & x(564) & x(565) & x(566) & x(567) & x(568) & x(569) & x(578) & x(580) & x(583) & x(584) & x(594) & x(597) & x(609) & x(610) & x(611) & x(620) & x(622) & x(624) & x(638) & x(665) & x(666) & x(668) & x(696) & x(697) & x(733) & x(737) & x(738) & x(740) & x(742) & x(767);
    y(96) <= not(p96_out);
    p96 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01111111111110100000000000111111111111111111111111111111111111111111111111111111",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 2,
            B => 139,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p96_in,
            y(0) => p96_out,
            y(1 to 14 - 1) => dummy96
        );


    p97_in <= x(247) & x(248) & x(249) & x(275) & x(276) & x(277) & x(278) & x(293) & x(294) & x(303) & x(304) & x(305) & x(306) & x(307) & x(320) & x(321) & x(322) & x(333) & x(334) & x(341) & x(342) & x(401) & x(403) & x(404) & x(454) & x(473) & x(501) & x(697) & x(718);
    y(97) <= not(p97_out);
    p97 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000000000011111110",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100101111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011000000010001010110010101110111111010000100010101100101011101111011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -90,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p97_in,
            y(0) => p97_out,
            y(1 to 14 - 1) => dummy97
        );


    p98_in <= x(44) & x(65) & x(94) & x(96) & x(97) & x(98) & x(102) & x(118) & x(121) & x(122) & x(123) & x(124) & x(125) & x(135) & x(147) & x(148) & x(171) & x(174) & x(238) & x(248) & x(266) & x(267) & x(276) & x(283) & x(291) & x(293) & x(294) & x(310) & x(321) & x(329) & x(330) & x(331) & x(332) & x(338) & x(346) & x(347) & x(348) & x(361) & x(366) & x(374) & x(375) & x(389) & x(390) & x(391) & x(396) & x(418) & x(446) & x(474) & x(475) & x(502) & x(524) & x(551) & x(619) & x(668) & x(705) & x(706) & x(707) & x(708) & x(744) & x(745) & x(746) & x(747) & x(750) & x(774);
    y(98) <= not(p98_out);
    p98 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000000000100000100101000000000111001100010000000000000000000",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101101011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101101110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 2,
            B => -202,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p98_in,
            y(0) => p98_out,
            y(1 to 14 - 1) => dummy98
        );


    p99_in <= x(92) & x(118) & x(120) & x(145) & x(192) & x(248) & x(249) & x(276) & x(277) & x(298) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(332) & x(333) & x(334) & x(357) & x(358) & x(359) & x(360) & x(386) & x(387) & x(388) & x(415) & x(425) & x(427) & x(454) & x(455) & x(468) & x(498) & x(514) & x(521) & x(612);
    y(99) <= not(p99_out);
    p99 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111100000100111110011111111111111111",
            TABLE => "000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 2,
            B => 51,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p99_in,
            y(0) => p99_out,
            y(1 to 13 - 1) => dummy99
        );


    p100_in <= x(127) & x(192) & x(198) & x(221) & x(248) & x(249) & x(276) & x(277) & x(296) & x(304) & x(305) & x(306) & x(317) & x(318) & x(319) & x(333) & x(338) & x(342) & x(343) & x(344) & x(345) & x(346) & x(347) & x(348) & x(366) & x(369) & x(370) & x(371) & x(372) & x(373) & x(375) & x(389) & x(390) & x(391) & x(396) & x(398) & x(399) & x(418) & x(446) & x(473) & x(474) & x(501) & x(517) & x(528) & x(529) & x(546) & x(557) & x(655) & x(656) & x(657) & x(681);
    y(100) <= not(p100_out);
    p100 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101000001000000010000000100000011100011111111110000",
            TABLE => "100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 2,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p100_in,
            y(0) => p100_out,
            y(1 to 13 - 1) => dummy100
        );


    p101_in <= x(35) & x(41) & x(46) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(77) & x(78) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(107) & x(108) & x(136) & x(171) & x(192) & x(199) & x(218) & x(220) & x(221) & x(248) & x(249) & x(273) & x(274) & x(275) & x(276) & x(277) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(332) & x(334) & x(350) & x(357) & x(358) & x(359) & x(360) & x(386) & x(387) & x(388) & x(415) & x(416) & x(443) & x(444) & x(446) & x(528) & x(543) & x(582) & x(607) & x(610) & x(611) & x(634) & x(636) & x(637) & x(638) & x(665) & x(697) & x(747);
    y(101) <= not(p101_out);
    p101 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000000000000101011111111111100000100000000000011011111111110",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111101110101001101010001000000110101000100000001000000000000001011110111010100110101000100001011010100010000100100001000101011011010011001011010010110011010011001011001101001011010011001011000010111000000010111111100010111000000010000000000010111000000010001011110000001011111100001011110000001111010000001011110000001100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000100000001000000011101000100000001110100011101000111111100001011110000001100000011110100010000001111010001110100001111110011010011001011010010110011010011001011001101001011010011001011011101000111111101000000011101000100000001110100000000000100000001110100001111110100000011110100010000001111010000001011110000001011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100110111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000010001010110010101110111111010000100010101100101011101111011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 2,
            B => -81,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p101_in,
            y(0) => p101_out,
            y(1 to 14 - 1) => dummy101
        );


    p102_in <= x(35) & x(46) & x(47) & x(69) & x(70) & x(72) & x(73) & x(74) & x(75) & x(78) & x(94) & x(95) & x(99) & x(101) & x(102) & x(152) & x(162) & x(163) & x(190) & x(191) & x(192) & x(218) & x(248) & x(276) & x(277) & x(305) & x(321) & x(322) & x(328) & x(329) & x(330) & x(331) & x(332) & x(354) & x(355) & x(357) & x(358) & x(359) & x(360) & x(387) & x(501) & x(513) & x(541) & x(542) & x(611) & x(697) & x(720) & x(740) & x(746);
    y(102) <= not(p102_out);
    p102 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111111111111111000000000011111111111111011100111",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 2,
            B => 74,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p102_in,
            y(0) => p102_out,
            y(1 to 13 - 1) => dummy102
        );


    p103_in <= x(333) & x(418) & x(426) & x(446) & x(453) & x(454) & x(501) & x(611) & x(658) & x(659) & x(686) & x(687) & x(688) & x(733);
    y(103) <= not(p103_out);
    p103 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01111111000001",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 3,
            B => 34,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p103_in,
            y(0) => p103_out,
            y(1 to 12 - 1) => dummy103
        );


    p104_in <= x(66) & x(244) & x(245) & x(271) & x(276) & x(277) & x(304) & x(305) & x(306) & x(330) & x(358) & x(367) & x(369) & x(406) & x(434) & x(493) & x(513);
    y(104) <= not(p104_out);
    p104 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111100110010",
            TABLE => "00000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000010000000100000011010100010000001101010011010100111111010010101101000010010000101101010001000010110101001101010010111101100101100110100101101001100101100110100110010110100101100110100110110010001000001111101110110010101100100010010011011011101100101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 78,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p104_in,
            y(0) => p104_out,
            y(1 to 14 - 1) => dummy104
        );


    p105_in <= x(35) & x(46) & x(47) & x(63) & x(64) & x(66) & x(68) & x(90) & x(91) & x(93) & x(105) & x(106) & x(130) & x(192) & x(220) & x(228) & x(229) & x(248) & x(256) & x(276) & x(277) & x(295) & x(304) & x(305) & x(306) & x(311) & x(323) & x(338) & x(341) & x(411) & x(446) & x(474) & x(501) & x(502) & x(526) & x(530) & x(540) & x(541) & x(542) & x(554) & x(558) & x(582) & x(608) & x(695) & x(718) & x(719) & x(720) & x(721) & x(722) & x(724) & x(748);
    y(105) <= not(p105_out);
    p105 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111111111001011011100010000010111101111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 3,
            B => 151,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p105_in,
            y(0) => p105_out,
            y(1 to 14 - 1) => dummy105
        );


    p106_in <= x(248) & x(274) & x(275) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(330) & x(333) & x(334) & x(358) & x(359) & x(390) & x(418) & x(439) & x(446) & x(528);
    y(106) <= not(p106_out);
    p106 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111110110011111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 4,
            B => 185,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p106_in,
            y(0) => p106_out,
            y(1 to 14 - 1) => dummy106
        );


    p107_in <= x(107) & x(249) & x(250) & x(276) & x(277) & x(294) & x(304) & x(305) & x(306) & x(316) & x(329) & x(330) & x(331) & x(333) & x(334) & x(343) & x(357) & x(358) & x(359) & x(360) & x(362) & x(369) & x(370) & x(387) & x(388) & x(390) & x(397) & x(398) & x(418) & x(425) & x(446) & x(451) & x(454) & x(455) & x(473) & x(474) & x(485) & x(501) & x(502) & x(529) & x(709) & x(710) & x(711) & x(712) & x(720) & x(721) & x(737) & x(745) & x(750);
    y(107) <= not(p107_out);
    p107 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000000001111001111101111011010011001000000000000",
            TABLE => "1110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101100111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010011000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 2,
            B => -62,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p107_in,
            y(0) => p107_out,
            y(1 to 13 - 1) => dummy107
        );


    p108_in <= x(98) & x(101) & x(102) & x(124) & x(125) & x(135) & x(152) & x(153) & x(192) & x(220) & x(221) & x(247) & x(248) & x(249) & x(275) & x(276) & x(277) & x(304) & x(305) & x(306) & x(315) & x(328) & x(329) & x(330) & x(331) & x(342) & x(343) & x(347) & x(357) & x(358) & x(359) & x(360) & x(370) & x(474) & x(502) & x(513) & x(720) & x(742);
    y(108) <= not(p108_out);
    p108 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000100111111111111100001110000100000",
            TABLE => "111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 3,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p108_in,
            y(0) => p108_out,
            y(1 to 14 - 1) => dummy108
        );


    p109_in <= x(44) & x(171) & x(178) & x(192) & x(221) & x(245) & x(247) & x(248) & x(249) & x(250) & x(274) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(321) & x(329) & x(330) & x(333) & x(334) & x(357) & x(358) & x(359) & x(360) & x(366) & x(387) & x(390) & x(418) & x(450) & x(451) & x(463) & x(469) & x(470) & x(479) & x(486) & x(487) & x(489) & x(490) & x(507) & x(508) & x(514) & x(515) & x(516) & x(517) & x(518) & x(525) & x(535) & x(536) & x(537) & x(564) & x(565) & x(592) & x(620) & x(629) & x(648) & x(649) & x(651) & x(675) & x(676) & x(677) & x(678) & x(704) & x(705) & x(706) & x(707) & x(709) & x(710) & x(724) & x(750);
    y(109) <= not(p109_out);
    p109 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000000000000000011001111010000100011110011111000000001000000000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 2,
            B => -187,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p109_in,
            y(0) => p109_out,
            y(1 to 14 - 1) => dummy109
        );


    p110_in <= x(207) & x(228) & x(247) & x(248) & x(267) & x(275) & x(276) & x(277) & x(295) & x(296) & x(305) & x(306) & x(311) & x(323) & x(359) & x(376) & x(390) & x(403) & x(418) & x(422) & x(441) & x(528) & x(554) & x(581) & x(582) & x(583) & x(609) & x(610) & x(611) & x(634) & x(638) & x(666) & x(676) & x(679) & x(697) & x(705) & x(706) & x(708) & x(709);
    y(110) <= not(p110_out);
    p110 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101101110011000111100111111111110010000",
            TABLE => "000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 3,
            B => 52,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p110_in,
            y(0) => p110_out,
            y(1 to 14 - 1) => dummy110
        );


    p111_in <= x(65) & x(106) & x(107) & x(248) & x(249) & x(276) & x(277) & x(294) & x(295) & x(304) & x(305) & x(306) & x(320) & x(321) & x(329) & x(330) & x(331) & x(332) & x(333) & x(334) & x(339) & x(357) & x(358) & x(359) & x(360) & x(366) & x(386) & x(387) & x(426) & x(427) & x(428) & x(430) & x(454) & x(455) & x(456) & x(457) & x(458) & x(483) & x(484) & x(485) & x(486) & x(487) & x(488) & x(513) & x(514) & x(515) & x(516) & x(543) & x(654) & x(665) & x(675) & x(676) & x(682) & x(685) & x(686) & x(704) & x(724);
    y(111) <= not(p111_out);
    p111 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000111111111110000111000010000000000000000000000101111111",
            TABLE => "011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => 1,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p111_in,
            y(0) => p111_out,
            y(1 to 12 - 1) => dummy111
        );


    p112_in <= x(35) & x(46) & x(50) & x(66) & x(91) & x(247) & x(248) & x(249) & x(275) & x(276) & x(277) & x(278) & x(293) & x(303) & x(304) & x(305) & x(306) & x(320) & x(321) & x(332) & x(333) & x(341) & x(387) & x(424) & x(446) & x(474) & x(489) & x(501) & x(502) & x(557) & x(558) & x(718) & x(719) & x(745);
    y(112) <= not(p112_out);
    p112 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000000000000000000011111111000",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011000000011101000100000011110100010010110011010010000000000000000",
            SHIFT => 3,
            B => -139,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p112_in,
            y(0) => p112_out,
            y(1 to 14 - 1) => dummy112
        );


    p113_in <= x(93) & x(145) & x(210) & x(211) & x(218) & x(233) & x(234) & x(256) & x(261) & x(322) & x(333) & x(350) & x(351) & x(354) & x(378) & x(379) & x(380) & x(382) & x(387) & x(388) & x(397) & x(406) & x(407) & x(416) & x(418) & x(433) & x(434) & x(435) & x(444) & x(446) & x(462) & x(472) & x(473) & x(487) & x(488) & x(500) & x(501) & x(514) & x(527) & x(528) & x(529) & x(583) & x(599) & x(611) & x(628) & x(629) & x(634) & x(659) & x(695) & x(697) & x(716) & x(718) & x(719) & x(720) & x(721) & x(740) & x(746);
    y(113) <= not(p113_out);
    p113 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011100000111111111000110011100100110010000000000101111111",
            TABLE => "000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => 2,
            B => -34,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p113_in,
            y(0) => p113_out,
            y(1 to 13 - 1) => dummy113
        );


    p114_in <= x(124) & x(146) & x(147) & x(159) & x(160) & x(238) & x(248) & x(249) & x(266) & x(267) & x(268) & x(269) & x(277) & x(295) & x(296) & x(306) & x(309) & x(310) & x(311) & x(316) & x(338) & x(345) & x(350) & x(356) & x(357) & x(358) & x(366) & x(376) & x(377) & x(389) & x(391) & x(418) & x(446) & x(473) & x(474) & x(501) & x(502) & x(528) & x(529) & x(557) & x(584) & x(612) & x(705) & x(736) & x(742) & x(743) & x(745) & x(746) & x(774);
    y(114) <= not(p114_out);
    p114 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001101100001001000101111101100000000000000000000",
            TABLE => "1011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010010000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 2,
            B => -110,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p114_in,
            y(0) => p114_out,
            y(1 to 13 - 1) => dummy114
        );


    p115_in <= x(239) & x(266) & x(267) & x(276) & x(277) & x(295) & x(304) & x(305) & x(342) & x(343) & x(358) & x(359) & x(360) & x(370) & x(387) & x(390) & x(418) & x(474) & x(502) & x(529) & x(557) & x(584) & x(666) & x(668) & x(733) & x(742);
    y(115) <= not(p115_out);
    p115 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111000000011111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 3,
            B => 69,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p115_in,
            y(0) => p115_out,
            y(1 to 13 - 1) => dummy115
        );


    p116_in <= x(171) & x(174) & x(178) & x(199) & x(242) & x(243) & x(244) & x(245) & x(249) & x(255) & x(256) & x(269) & x(270) & x(271) & x(272) & x(273) & x(274) & x(277) & x(283) & x(296) & x(297) & x(300) & x(301) & x(304) & x(305) & x(306) & x(309) & x(310) & x(311) & x(312) & x(333) & x(338) & x(339) & x(357) & x(358) & x(359) & x(360) & x(362) & x(366) & x(387) & x(390) & x(403) & x(405) & x(406) & x(407) & x(418) & x(433) & x(434) & x(446) & x(459) & x(474) & x(479) & x(481) & x(486) & x(507) & x(515) & x(516) & x(535) & x(625) & x(676) & x(677) & x(678) & x(679) & x(692) & x(695) & x(704) & x(705) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(774);
    y(116) <= not(p116_out);
    p116 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000000000000000000000011110010111101101000101100000011000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 2,
            B => -124,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p116_in,
            y(0) => p116_out,
            y(1 to 14 - 1) => dummy116
        );


    p117_in <= x(66) & x(105) & x(106) & x(192) & x(228) & x(242) & x(249) & x(255) & x(256) & x(268) & x(269) & x(270) & x(276) & x(277) & x(297) & x(298) & x(299) & x(300) & x(302) & x(305) & x(310) & x(311) & x(330) & x(331) & x(332) & x(338) & x(358) & x(359) & x(360) & x(361) & x(366) & x(387) & x(388) & x(389) & x(407) & x(431) & x(446) & x(475) & x(720) & x(774);
    y(117) <= not(p117_out);
    p117 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111001000001100000100000000000000110010",
            TABLE => "0000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010011011001000100000101100100010010010010110011010010000000000000000",
            SHIFT => 3,
            B => -72,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p117_in,
            y(0) => p117_out,
            y(1 to 14 - 1) => dummy117
        );


    p118_in <= x(218) & x(228) & x(251) & x(277) & x(278) & x(306) & x(310) & x(311) & x(316) & x(322) & x(338) & x(343) & x(350) & x(351) & x(352) & x(366) & x(378) & x(379) & x(389) & x(391) & x(399) & x(407) & x(416) & x(418) & x(425) & x(426) & x(428) & x(444) & x(446) & x(453) & x(454) & x(473) & x(474) & x(482) & x(501) & x(502) & x(528) & x(529) & x(557) & x(691) & x(695) & x(697) & x(719) & x(720);
    y(118) <= not(p118_out);
    p118 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00111100110111101100010000000000000000011011",
            TABLE => "000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 2,
            B => -80,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p118_in,
            y(0) => p118_out,
            y(1 to 13 - 1) => dummy118
        );


    p119_in <= x(35) & x(62) & x(63) & x(64) & x(65) & x(66) & x(68) & x(106) & x(107) & x(108) & x(135) & x(145) & x(147) & x(171) & x(184) & x(201) & x(211) & x(212) & x(228) & x(229) & x(256) & x(269) & x(270) & x(271) & x(272) & x(276) & x(283) & x(297) & x(298) & x(299) & x(301) & x(311) & x(339) & x(361) & x(409) & x(422) & x(424) & x(437) & x(445) & x(465) & x(501) & x(535) & x(666) & x(668) & x(677) & x(679) & x(695) & x(732) & x(738) & x(740);
    y(119) <= not(p119_out);
    p119 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111111000101100000001000000000000101011001111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 2,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p119_in,
            y(0) => p119_out,
            y(1 to 13 - 1) => dummy119
        );


    p120_in <= x(95) & x(96) & x(98) & x(163) & x(191) & x(192) & x(221) & x(222) & x(248) & x(249) & x(303) & x(329) & x(330) & x(331) & x(332) & x(358) & x(359) & x(611) & x(705) & x(707) & x(717) & x(718) & x(719) & x(720) & x(721) & x(741) & x(742) & x(744) & x(745) & x(746) & x(747);
    y(120) <= not(p120_out);
    p120 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001111111000000010000000000000",
            TABLE => "0111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => -131,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p120_in,
            y(0) => p120_out,
            y(1 to 14 - 1) => dummy120
        );


    p121_in <= x(95) & x(108) & x(211) & x(248) & x(249) & x(250) & x(256) & x(277) & x(278) & x(305) & x(322) & x(350) & x(351) & x(354) & x(359) & x(360) & x(379) & x(387) & x(388) & x(389) & x(397) & x(399) & x(415) & x(416) & x(417) & x(418) & x(425) & x(426) & x(427) & x(443) & x(444) & x(446) & x(453) & x(454) & x(471) & x(472) & x(473) & x(481) & x(482) & x(488) & x(501) & x(508) & x(509) & x(510) & x(511) & x(527) & x(528) & x(529) & x(538) & x(539) & x(545) & x(546) & x(553) & x(554) & x(557) & x(564) & x(567) & x(568) & x(581) & x(583) & x(695) & x(697) & x(719) & x(720) & x(722);
    y(121) <= not(p121_out);
    p121 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00111101111111001000000000000000000000010000000000000000000010111",
            TABLE => "00010111011111110000000100010111000000010001011100000000000000010001011101111110100000010001011110000001000101111110100010000001100101100110100101101001100101100110100110010110100101100110100100000001000101110001011101111111000000000000000100000001000101111000000100010111000101110111111011101000100000011000000100010111011010011001011010010110011010011001011001101001011010011001011000100000000000001011001000100000101100100010000011111011101100100010010001001101101100100010010010110010001001001101101110110010011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111101111100011101000111000001000100011100000100000001000000000001110011110001110100011100001100010001110000110000001100001110001011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100010111000000010111111100010111000101111000000101111110000101111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 2,
            B => -88,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p121_in,
            y(0) => p121_out,
            y(1 to 14 - 1) => dummy121
        );


    p122_in <= x(35) & x(63) & x(64) & x(66) & x(68) & x(91) & x(92) & x(172) & x(276) & x(277) & x(304) & x(305) & x(324) & x(330) & x(352) & x(387) & x(411) & x(415) & x(416) & x(526) & x(554) & x(581) & x(606) & x(607) & x(632) & x(634) & x(636) & x(647) & x(659) & x(685) & x(686) & x(724) & x(767);
    y(122) <= not(p122_out);
    p122 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000010000111010000000000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 3,
            B => -152,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p122_in,
            y(0) => p122_out,
            y(1 to 14 - 1) => dummy122
        );


    p123_in <= x(249) & x(277) & x(305) & x(329) & x(330) & x(331) & x(342) & x(357) & x(358) & x(359) & x(360) & x(369) & x(370) & x(387) & x(473) & x(474) & x(489) & x(501) & x(516) & x(529) & x(611);
    y(123) <= not(p123_out);
    p123 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111000000000001111111",
            TABLE => "000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 3,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p123_in,
            y(0) => p123_out,
            y(1 to 13 - 1) => dummy123
        );


    p124_in <= x(44) & x(145) & x(178) & x(203) & x(205) & x(206) & x(207) & x(234) & x(243) & x(247) & x(248) & x(276) & x(277) & x(303) & x(304) & x(305) & x(306) & x(310) & x(314) & x(315) & x(333) & x(334) & x(338) & x(339) & x(342) & x(357) & x(358) & x(359) & x(360) & x(362) & x(366) & x(378) & x(379) & x(390) & x(391) & x(408) & x(418) & x(489) & x(490) & x(521) & x(582) & x(695) & x(704) & x(724) & x(764) & x(774);
    y(124) <= not(p124_out);
    p124 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100000000000000000000000111100110010110010000",
            TABLE => "1110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010010100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101101110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 3,
            B => -134,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p124_in,
            y(0) => p124_out,
            y(1 to 14 - 1) => dummy124
        );


    p125_in <= x(181) & x(182) & x(211) & x(212) & x(229) & x(248) & x(249) & x(250) & x(276) & x(277) & x(303) & x(304) & x(305) & x(306) & x(322) & x(332) & x(333) & x(334) & x(350) & x(359) & x(362) & x(377) & x(387) & x(397) & x(399) & x(547) & x(695) & x(705) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(732) & x(744) & x(745) & x(746) & x(747) & x(748) & x(750);
    y(125) <= not(p125_out);
    p125 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000010000000000000010011110000000000000000",
            TABLE => "111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => -163,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p125_in,
            y(0) => p125_out,
            y(1 to 14 - 1) => dummy125
        );


    p126_in <= x(73) & x(91) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(118) & x(136) & x(191) & x(192) & x(202) & x(220) & x(221) & x(228) & x(248) & x(249) & x(256) & x(275) & x(276) & x(277) & x(294) & x(295) & x(296) & x(304) & x(305) & x(306) & x(310) & x(316) & x(328) & x(329) & x(330) & x(331) & x(334) & x(338) & x(339) & x(343) & x(344) & x(366) & x(375) & x(383) & x(384) & x(385) & x(398) & x(401) & x(418) & x(428) & x(474) & x(501) & x(529) & x(544) & x(705) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(774);
    y(126) <= not(p126_out);
    p126 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000001110110110111000111010000100110111111010000000000000",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100100000100010011010000000000000100010011011101111100000100010011010010010001001101101100100010010001001101110110110010010001001101100101100110100101101001100101100110100110010110100101100110100101000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011000001000000000001000111000001000100011100000100011101111100011100001100001110001100011100001100010001110000110001110011110001110011010011001011010010110011010011001011001101001011010011001011011010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100100000001000101110000000000000001000101110111111100000001000101111000000100010111111010001000000100010111011111101000000100010111011010011001011010010110011010011001011001101001011010011001011000001000000000001000111000001000100011100000100011101111100011100001100001110001100011100001100010001110000110001110011110001110011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 2,
            B => -98,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p126_in,
            y(0) => p126_out,
            y(1 to 14 - 1) => dummy126
        );


    p127_in <= x(64) & x(66) & x(144) & x(276) & x(277) & x(303) & x(306) & x(310) & x(331) & x(338) & x(343) & x(358) & x(359) & x(360) & x(366) & x(386) & x(387) & x(388) & x(415) & x(416) & x(418) & x(444) & x(694) & x(695) & x(720);
    y(127) <= not(p127_out);
    p127 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101111111111111111111000",
            TABLE => "0000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => 130,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p127_in,
            y(0) => p127_out,
            y(1 to 13 - 1) => dummy127
        );


    p128_in <= x(108) & x(145) & x(152) & x(154) & x(198) & x(235) & x(248) & x(250) & x(262) & x(263) & x(264) & x(277) & x(290) & x(306) & x(321) & x(322) & x(326) & x(338) & x(348) & x(349) & x(350) & x(366) & x(417) & x(473) & x(474) & x(501) & x(529) & x(546) & x(547) & x(573) & x(574) & x(575) & x(600) & x(601) & x(602) & x(650) & x(660) & x(661) & x(662) & x(666);
    y(128) <= not(p128_out);
    p128 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000110011101000010001111111111111100001",
            TABLE => "0111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101100010101110111111000000100010101100000010001010110000000000000010001010111011110101000010001010110100001000101011110101000100001001101001100101101001011001101001100101100110100101101001100101101101010001000000010000000000000011111101110101001101010001000000110101000100001001000010001010111011110111010100110101000100001010010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101101010001000000110101000100001010010110011010010000000000000000",
            SHIFT => 2,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p128_in,
            y(0) => p128_out,
            y(1 to 13 - 1) => dummy128
        );


    p129_in <= x(165) & x(182) & x(183) & x(184) & x(192) & x(193) & x(198) & x(210) & x(211) & x(221) & x(248) & x(249) & x(250) & x(263) & x(264) & x(276) & x(277) & x(278) & x(292) & x(303) & x(304) & x(305) & x(306) & x(310) & x(332) & x(333) & x(334) & x(338) & x(349) & x(350) & x(366) & x(377) & x(378) & x(405) & x(406) & x(411) & x(418) & x(438) & x(446) & x(465) & x(473) & x(474) & x(501) & x(510) & x(537) & x(774);
    y(129) <= not(p129_out);
    p129 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111110111111001110111101110110111100000000110",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010010000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 2,
            B => 29,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p129_in,
            y(0) => p129_out,
            y(1 to 13 - 1) => dummy129
        );


    p130_in <= x(319) & x(330) & x(331) & x(332) & x(338) & x(345) & x(346) & x(347) & x(357) & x(358) & x(359) & x(360) & x(371) & x(372) & x(373) & x(387) & x(399) & x(400) & x(414) & x(442) & x(443) & x(471) & x(473) & x(497) & x(498) & x(501) & x(529) & x(584) & x(611) & x(638) & x(666);
    y(130) <= not(p130_out);
    p130 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000100000000000000000100111111",
            TABLE => "1111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 2,
            B => -36,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p130_in,
            y(0) => p130_out,
            y(1 to 13 - 1) => dummy130
        );


    p131_in <= x(65) & x(71) & x(90) & x(136) & x(165) & x(182) & x(183) & x(203) & x(210) & x(211) & x(221) & x(228) & x(229) & x(249) & x(250) & x(256) & x(276) & x(277) & x(297) & x(299) & x(304) & x(305) & x(306) & x(310) & x(311) & x(333) & x(334) & x(338) & x(339) & x(343) & x(350) & x(359) & x(360) & x(362) & x(366) & x(369) & x(370) & x(378) & x(387) & x(388) & x(390) & x(396) & x(397) & x(405) & x(416) & x(418) & x(451) & x(466) & x(479) & x(695) & x(704) & x(717) & x(720) & x(721);
    y(131) <= not(p131_out);
    p131 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111101110011011001110011000100100010010010110110111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 2,
            B => 16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p131_in,
            y(0) => p131_out,
            y(1 to 13 - 1) => dummy131
        );


    p132_in <= x(66) & x(276) & x(277) & x(304) & x(305) & x(306) & x(329) & x(330) & x(331) & x(332) & x(355) & x(356) & x(357) & x(358) & x(359) & x(360) & x(484) & x(528) & x(704) & x(705) & x(712) & x(718) & x(724) & x(747);
    y(132) <= not(p132_out);
    p132 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111000000000001111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => 34,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p132_in,
            y(0) => p132_out,
            y(1 to 13 - 1) => dummy132
        );


    p133_in <= x(108) & x(165) & x(192) & x(219) & x(220) & x(245) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(278) & x(305) & x(306) & x(328) & x(329) & x(333) & x(334) & x(338) & x(358) & x(359) & x(360) & x(362) & x(366) & x(387) & x(388) & x(390) & x(418) & x(434) & x(507) & x(695);
    y(133) <= not(p133_out);
    p133 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011111111111111100111000110011000",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 3,
            B => 147,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p133_in,
            y(0) => p133_out,
            y(1 to 14 - 1) => dummy133
        );


    p134_in <= x(46) & x(63) & x(64) & x(66) & x(68) & x(90) & x(91) & x(144) & x(192) & x(199) & x(220) & x(221) & x(228) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(298) & x(302) & x(304) & x(305) & x(306) & x(309) & x(310) & x(311) & x(328) & x(329) & x(330) & x(331) & x(338) & x(357) & x(358) & x(359) & x(360) & x(366) & x(424) & x(445) & x(514) & x(546) & x(558) & x(628) & x(632) & x(634) & x(647) & x(664) & x(666) & x(683) & x(685) & x(696) & x(724) & x(767);
    y(134) <= not(p134_out);
    p134 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000001010010000001100011111111111111011100000000000",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100110001110000010001110111110001110000010000000000010001110000010001000111000011000111001111000111000011000011100011000111000011000100101100110100101101001100101100110100110010110100101100110100111101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011010000000111010001110100011111110000000001000000010000000111010001000000111101000111010000111111000010111100000011000000111101000100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000001000000000001011100000001000101110000000101111111000101111000000111101000000101111000000100010111100000010111111000010111011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -68,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p134_in,
            y(0) => p134_out,
            y(1 to 14 - 1) => dummy134
        );


    p135_in <= x(35) & x(38) & x(46) & x(63) & x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(78) & x(91) & x(93) & x(94) & x(95) & x(97) & x(106) & x(107) & x(108) & x(190) & x(192) & x(201) & x(210) & x(211) & x(218) & x(219) & x(220) & x(221) & x(244) & x(246) & x(247) & x(248) & x(249) & x(272) & x(273) & x(274) & x(275) & x(276) & x(277) & x(304) & x(305) & x(306) & x(320) & x(329) & x(333) & x(334) & x(347) & x(348) & x(358) & x(359) & x(360) & x(369) & x(387) & x(388) & x(396) & x(397) & x(424) & x(445) & x(473) & x(487) & x(501) & x(514) & x(515) & x(516) & x(543) & x(544) & x(675) & x(742) & x(746);
    y(135) <= not(p135_out);
    p135 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111111111111111100011000000000000000000010000111011000111111111011",
            TABLE => "00000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000100000001000000011101000100000001110100011101000111111100001011110000001100000011110100010000001111010001110100001111110011010011001011010010110011010011001011001101001011010011001011010000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111101111100011101000111000001000100011100000100000001000000000001110011110001110100011100001100010001110000110000001100001110001011010011001011010010110011010011001011001101001011010011001011000101011101111110000001000101011000000100010101100000000000000100010101110111101010000100010101101000010001010111101010001000010011010011001011010010110011010011001011001101001011010011001011001000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100010000011100010111000111110111000110000111000101110001111001111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 2,
            B => 27,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p135_in,
            y(0) => p135_out,
            y(1 to 14 - 1) => dummy135
        );


    p136_in <= x(106) & x(145) & x(220) & x(237) & x(238) & x(247) & x(248) & x(276) & x(277) & x(302) & x(305) & x(328) & x(329) & x(330) & x(331) & x(332) & x(350) & x(357) & x(358) & x(359) & x(360) & x(361) & x(389) & x(390) & x(418) & x(446) & x(452) & x(474) & x(475) & x(479) & x(480) & x(502) & x(507) & x(558) & x(619) & x(622);
    y(136) <= not(p136_out);
    p136 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010110000101111111111111111111111111",
            TABLE => "001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => 123,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p136_in,
            y(0) => p136_out,
            y(1 to 14 - 1) => dummy136
        );


    p137_in <= x(249) & x(250) & x(277) & x(278) & x(305) & x(306) & x(309) & x(329) & x(330) & x(333) & x(349) & x(350) & x(357) & x(358) & x(359) & x(386) & x(387) & x(388) & x(404) & x(406) & x(407) & x(412) & x(414) & x(415) & x(426) & x(433) & x(435) & x(441) & x(454) & x(455) & x(482) & x(501) & x(507) & x(529) & x(612) & x(647) & x(688);
    y(137) <= not(p137_out);
    p137 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111110001110000001110000110000010011",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101101000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010011101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 2,
            B => -28,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p137_in,
            y(0) => p137_out,
            y(1 to 13 - 1) => dummy137
        );


    p138_in <= x(93) & x(220) & x(221) & x(248) & x(249) & x(250) & x(256) & x(276) & x(277) & x(278) & x(304) & x(305) & x(306) & x(310) & x(328) & x(329) & x(330) & x(331) & x(333) & x(334) & x(338) & x(357) & x(358) & x(359) & x(360) & x(366) & x(387) & x(388) & x(453) & x(454) & x(501) & x(613) & x(675) & x(742);
    y(138) <= not(p138_out);
    p138 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111110111111000001100000000000010",
            TABLE => "0000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101101110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011011001000100000101100100010010010010110011010010000000000000000",
            SHIFT => 3,
            B => -41,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p138_in,
            y(0) => p138_out,
            y(1 to 14 - 1) => dummy138
        );


    p139_in <= x(39) & x(180) & x(181) & x(182) & x(184) & x(185) & x(200) & x(208) & x(228) & x(247) & x(248) & x(256) & x(275) & x(276) & x(277) & x(304) & x(305) & x(311) & x(360) & x(361) & x(388) & x(463) & x(474) & x(619) & x(719) & x(721) & x(723) & x(732) & x(733);
    y(139) <= not(p139_out);
    p139 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111101011011111000000011111",
            TABLE => "00000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100101011000000101011111100101011000000100000000000101011000000100010101101000010101111010010101101000010110101000010101101000010011010011001011010010110011010011001011001101001011010011001011000000000000000100000001000101011000000100010101100101011101111111101010001000010010000100010101101000010001010110010101110111101011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100000001000101110001011101111111100000010001011100010111011111100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 3,
            B => 17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p139_in,
            y(0) => p139_out,
            y(1 to 14 - 1) => dummy139
        );


    p140_in <= x(35) & x(40) & x(64) & x(66) & x(70) & x(97) & x(107) & x(108) & x(136) & x(192) & x(214) & x(215) & x(216) & x(217) & x(218) & x(220) & x(221) & x(242) & x(243) & x(244) & x(245) & x(246) & x(248) & x(249) & x(273) & x(274) & x(276) & x(277) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(332) & x(334) & x(357) & x(358) & x(359) & x(360) & x(386) & x(387) & x(388) & x(445) & x(509) & x(510) & x(514) & x(515) & x(542) & x(543) & x(596) & x(675) & x(676) & x(704) & x(746);
    y(140) <= not(p140_out);
    p140 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000011111111111111111111110000010000000011000011110",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 2,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p140_in,
            y(0) => p140_out,
            y(1 to 13 - 1) => dummy140
        );


    p141_in <= x(72) & x(171) & x(213) & x(242) & x(267) & x(292) & x(368) & x(369) & x(370) & x(397) & x(398) & x(406) & x(414) & x(415) & x(434) & x(442) & x(443) & x(453) & x(473) & x(535) & x(705) & x(732) & x(733) & x(735) & x(736) & x(742) & x(746);
    y(141) <= not(p141_out);
    p141 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011110111110110111011111111",
            TABLE => "000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => 3,
            B => 108,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p141_in,
            y(0) => p141_out,
            y(1 to 13 - 1) => dummy141
        );


    p142_in <= x(35) & x(40) & x(46) & x(64) & x(66) & x(74) & x(276) & x(303) & x(331) & x(332) & x(359) & x(360) & x(387) & x(388) & x(415) & x(416) & x(443) & x(444) & x(475) & x(489) & x(490) & x(491) & x(500) & x(518) & x(558) & x(584) & x(611) & x(629) & x(666) & x(682) & x(686) & x(742);
    y(142) <= not(p142_out);
    p142 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000000011110111101001",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 3,
            B => -76,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p142_in,
            y(0) => p142_out,
            y(1 to 14 - 1) => dummy142
        );


    p143_in <= x(109) & x(157) & x(190) & x(192) & x(248) & x(249) & x(276) & x(277) & x(304) & x(305) & x(306) & x(329) & x(330) & x(331) & x(358) & x(359) & x(360) & x(380) & x(463) & x(528) & x(569) & x(608);
    y(143) <= not(p143_out);
    p143 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000000011111111000",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011000000011101000100000011110100010010110011010010000000000000000",
            SHIFT => 3,
            B => -69,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p143_in,
            y(0) => p143_out,
            y(1 to 13 - 1) => dummy143
        );


    p144_in <= x(303) & x(304) & x(330) & x(331) & x(332) & x(341) & x(342) & x(369) & x(406) & x(473) & x(501) & x(516) & x(529) & x(611) & x(706) & x(707) & x(719) & x(745) & x(746);
    y(144) <= not(p144_out);
    p144 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111111100000011111",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => 67,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p144_in,
            y(0) => p144_out,
            y(1 to 13 - 1) => dummy144
        );


    p145_in <= x(79) & x(91) & x(108) & x(136) & x(203) & x(210) & x(211) & x(212) & x(216) & x(231) & x(232) & x(233) & x(276) & x(323) & x(350) & x(351) & x(378) & x(406) & x(444) & x(473) & x(489) & x(501) & x(528) & x(529) & x(575) & x(604) & x(695);
    y(145) <= not(p145_out);
    p145 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000101111000011111001000001",
            TABLE => "110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110110101001001011011111111",
            SHIFT => 2,
            B => -35,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p145_in,
            y(0) => p145_out,
            y(1 to 12 - 1) => dummy145
        );


    p146_in <= x(116) & x(220) & x(238) & x(248) & x(249) & x(276) & x(277) & x(306) & x(342) & x(343) & x(359) & x(369) & x(370) & x(371) & x(386) & x(387) & x(390) & x(391) & x(397) & x(398) & x(414) & x(415) & x(416) & x(418) & x(442) & x(443) & x(446) & x(474) & x(475) & x(502) & x(531) & x(557) & x(558) & x(613) & x(666) & x(697) & x(746);
    y(146) <= not(p146_out);
    p146 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010000000000000110000010011111111111",
            TABLE => "1110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 2,
            B => -29,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p146_in,
            y(0) => p146_out,
            y(1 to 13 - 1) => dummy146
        );


    p147_in <= x(64) & x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(91) & x(93) & x(94) & x(97) & x(106) & x(108) & x(136) & x(190) & x(192) & x(198) & x(220) & x(221) & x(248) & x(249) & x(276) & x(277) & x(278) & x(304) & x(305) & x(306) & x(331) & x(333) & x(334) & x(346) & x(347) & x(348) & x(349) & x(359) & x(360) & x(369) & x(370) & x(371) & x(375) & x(387) & x(388) & x(389) & x(396) & x(417) & x(418) & x(445) & x(473) & x(474) & x(501) & x(514) & x(515) & x(516) & x(517) & x(528) & x(529) & x(543) & x(544) & x(545) & x(546) & x(574) & x(613) & x(675) & x(676) & x(697) & x(738) & x(739) & x(742) & x(745);
    y(147) <= not(p147_out);
    p147 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111111100010000000000100000011000011101111111111111111110011111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 2,
            B => 63,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p147_in,
            y(0) => p147_out,
            y(1 to 14 - 1) => dummy147
        );


    p148_in <= x(151) & x(181) & x(186) & x(228) & x(229) & x(230) & x(248) & x(249) & x(256) & x(257) & x(258) & x(276) & x(277) & x(283) & x(284) & x(285) & x(304) & x(305) & x(310) & x(311) & x(312) & x(313) & x(330) & x(331) & x(338) & x(339) & x(358) & x(359) & x(360) & x(366) & x(376) & x(387) & x(388) & x(431) & x(694) & x(695) & x(720) & x(721) & x(732) & x(733) & x(769) & x(773) & x(774);
    y(148) <= not(p148_out);
    p148 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001110011100111001111111111110110000000111",
            TABLE => "0111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100010101110111111000000100010101100000010001010110000000000000010001010111011110101000010001010110100001000101011110101000100001001101001100101101001011001101001100101100110100101101001100101100000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010011111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => 82,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p148_in,
            y(0) => p148_out,
            y(1 to 14 - 1) => dummy148
        );


    p149_in <= x(35) & x(40) & x(63) & x(64) & x(66) & x(76) & x(78) & x(91) & x(107) & x(108) & x(235) & x(248) & x(249) & x(276) & x(277) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(333) & x(334) & x(338) & x(341) & x(343) & x(344) & x(357) & x(358) & x(359) & x(360) & x(366) & x(386) & x(387) & x(388) & x(414) & x(415) & x(416) & x(440) & x(441) & x(443) & x(444) & x(572) & x(601) & x(602) & x(705) & x(707) & x(738) & x(741) & x(742) & x(743) & x(745) & x(746) & x(774);
    y(149) <= not(p149_out);
    p149 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111110000001111001111111111111111111111111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 2,
            B => 126,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p149_in,
            y(0) => p149_out,
            y(1 to 13 - 1) => dummy149
        );


    p150_in <= x(98) & x(203) & x(233) & x(248) & x(276) & x(315) & x(330) & x(332) & x(338) & x(339) & x(342) & x(343) & x(350) & x(356) & x(366) & x(369) & x(370) & x(371) & x(378) & x(390) & x(396) & x(397) & x(398) & x(405) & x(418) & x(433) & x(466) & x(474) & x(479) & x(502) & x(573) & x(678) & x(720) & x(721);
    y(150) <= not(p150_out);
    p150 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111110011110011110011100010000100",
            TABLE => "0000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010010101110111111000000100010101100000010001010110000000000000010001010111011110101000010001010110100001000101011110101000100001001101001100101101001011001101001100101100110100101101001100101101110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101101000111000001000100011100001100010010110011010010000000000000000",
            SHIFT => 3,
            B => 38,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p150_in,
            y(0) => p150_out,
            y(1 to 14 - 1) => dummy150
        );


    p151_in <= x(65) & x(66) & x(67) & x(68) & x(69) & x(70) & x(71) & x(93) & x(106) & x(136) & x(192) & x(193) & x(198) & x(220) & x(221) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(304) & x(305) & x(306) & x(328) & x(329) & x(330) & x(333) & x(334) & x(338) & x(356) & x(357) & x(358) & x(359) & x(360) & x(366) & x(387) & x(388) & x(417) & x(445) & x(450) & x(473) & x(501) & x(510) & x(537) & x(742);
    y(151) <= not(p151_out);
    p151 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000001110111111111110001100000000000100110",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 3,
            B => -51,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p151_in,
            y(0) => p151_out,
            y(1 to 14 - 1) => dummy151
        );


    p152_in <= x(41) & x(46) & x(64) & x(66) & x(68) & x(69) & x(70) & x(90) & x(91) & x(99) & x(101) & x(103) & x(104) & x(162) & x(192) & x(208) & x(220) & x(221) & x(248) & x(249) & x(250) & x(276) & x(277) & x(304) & x(305) & x(306) & x(310) & x(320) & x(321) & x(322) & x(328) & x(330) & x(331) & x(332) & x(338) & x(339) & x(342) & x(358) & x(359) & x(360) & x(366) & x(368) & x(389) & x(390) & x(418) & x(424) & x(425) & x(440) & x(446) & x(453) & x(454) & x(474) & x(475) & x(484) & x(485) & x(502) & x(535) & x(620) & x(648) & x(649) & x(651) & x(675) & x(677) & x(704) & x(707) & x(709) & x(711) & x(712) & x(715) & x(722) & x(750);
    y(152) <= not(p152_out);
    p152 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000000000000000000011110001110011111011111111000000000000000",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100100001000100011101000111011101111000000000000100000001000100011100001100010001110100011101110011101110001000110000001100010001110011010011001011010010110011010011001011001101001011010011001011000000000000000100000001000101011000000100010101100101011101111111101010001000010010000100010101101000010001010110010101110111101011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100110000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -192,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p152_in,
            y(0) => p152_out,
            y(1 to 15 - 1) => dummy152
        );


    p153_in <= x(40) & x(46) & x(47) & x(48) & x(64) & x(66) & x(68) & x(74) & x(78) & x(105) & x(106) & x(145) & x(171) & x(172) & x(200) & x(201) & x(202) & x(211) & x(220) & x(228) & x(248) & x(256) & x(269) & x(270) & x(276) & x(277) & x(278) & x(283) & x(295) & x(296) & x(298) & x(299) & x(301) & x(302) & x(306) & x(310) & x(311) & x(326) & x(328) & x(338) & x(339) & x(366) & x(377) & x(403) & x(407) & x(424) & x(425) & x(426) & x(452) & x(453) & x(475) & x(480) & x(502) & x(507) & x(535) & x(558) & x(563) & x(564) & x(592) & x(619) & x(676) & x(677) & x(695) & x(705) & x(708) & x(772) & x(773) & x(774);
    y(153) <= not(p153_out);
    p153 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000111111001011100011111110111111100011111111111111111011111",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 2,
            B => 98,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p153_in,
            y(0) => p153_out,
            y(1 to 14 - 1) => dummy153
        );


    p154_in <= x(64) & x(66) & x(192) & x(220) & x(228) & x(247) & x(248) & x(249) & x(256) & x(275) & x(276) & x(277) & x(299) & x(303) & x(304) & x(305) & x(306) & x(328) & x(329) & x(330) & x(343) & x(350) & x(360) & x(361) & x(389) & x(502) & x(584) & x(666) & x(695) & x(717) & x(718) & x(719) & x(720) & x(721);
    y(154) <= not(p154_out);
    p154 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111011101110111100011000011111111",
            TABLE => "0000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010011000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 4,
            B => 185,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p154_in,
            y(0) => p154_out,
            y(1 to 15 - 1) => dummy154
        );


    p155_in <= x(48) & x(66) & x(276) & x(277) & x(293) & x(294) & x(305) & x(321) & x(322) & x(330) & x(331) & x(342) & x(350) & x(358) & x(360) & x(446) & x(473) & x(501) & x(528) & x(709) & x(719) & x(720) & x(721) & x(742) & x(745) & x(746) & x(747);
    y(155) <= not(p155_out);
    p155 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000000110011111100000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 3,
            B => -54,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p155_in,
            y(0) => p155_out,
            y(1 to 13 - 1) => dummy155
        );


    p156_in <= x(108) & x(292) & x(338) & x(361) & x(366) & x(391) & x(398) & x(399) & x(400) & x(415) & x(426) & x(427) & x(428) & x(470) & x(606) & x(694) & x(732);
    y(156) <= not(p156_out);
    p156 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01111100000000000",
            TABLE => "00000001000101110001011101111111000000000000000100000001000101111000000100010111000101110111111011101000100000011000000100010111011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -33,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p156_in,
            y(0) => p156_out,
            y(1 to 13 - 1) => dummy156
        );


    p157_in <= x(78) & x(106) & x(109) & x(171) & x(267) & x(294) & x(295) & x(296) & x(305) & x(310) & x(311) & x(332) & x(339) & x(354) & x(355) & x(358) & x(359) & x(360) & x(366) & x(418) & x(439) & x(446) & x(459) & x(467) & x(469) & x(473) & x(474) & x(501) & x(502) & x(528) & x(529) & x(557) & x(564) & x(592) & x(704) & x(708);
    y(157) <= not(p157_out);
    p157 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110000000001011111000010000000000000",
            TABLE => "100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => -119,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p157_in,
            y(0) => p157_out,
            y(1 to 14 - 1) => dummy157
        );


    p158_in <= x(165) & x(192) & x(193) & x(248) & x(249) & x(276) & x(277) & x(303) & x(304) & x(305) & x(306) & x(319) & x(333) & x(341) & x(342) & x(369) & x(418) & x(446) & x(473) & x(474) & x(475) & x(490) & x(501) & x(502) & x(518) & x(528) & x(529) & x(545) & x(546) & x(547) & x(574) & x(611) & x(695) & x(697) & x(705) & x(706) & x(707) & x(708) & x(709) & x(711) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(747) & x(750);
    y(158) <= not(p158_out);
    p158 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111111111100000000000000001011111111111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 3,
            B => 127,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p158_in,
            y(0) => p158_out,
            y(1 to 14 - 1) => dummy158
        );


    p159_in <= x(66) & x(135) & x(192) & x(220) & x(221) & x(248) & x(249) & x(276) & x(277) & x(278) & x(304) & x(305) & x(306) & x(321) & x(322) & x(328) & x(329) & x(330) & x(331) & x(333) & x(334) & x(339) & x(357) & x(358) & x(359) & x(360) & x(366) & x(389) & x(390) & x(418) & x(424) & x(425) & x(453) & x(454) & x(474) & x(475) & x(502) & x(668) & x(733);
    y(159) <= not(p159_out);
    p159 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111111111000011100001000000000000",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 3,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p159_in,
            y(0) => p159_out,
            y(1 to 14 - 1) => dummy159
        );


    p160_in <= x(75) & x(153) & x(154) & x(155) & x(161) & x(183) & x(198) & x(220) & x(235) & x(248) & x(249) & x(256) & x(276) & x(277) & x(305) & x(310) & x(312) & x(328) & x(329) & x(330) & x(331) & x(332) & x(338) & x(339) & x(357) & x(358) & x(359) & x(360) & x(366) & x(418) & x(438) & x(439) & x(473) & x(501) & x(513) & x(528);
    y(160) <= not(p160_out);
    p160 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111101000000000001111100111100000010",
            TABLE => "000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => -65,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p160_in,
            y(0) => p160_out,
            y(1 to 14 - 1) => dummy160
        );


    p161_in <= x(39) & x(93) & x(117) & x(118) & x(133) & x(135) & x(145) & x(147) & x(161) & x(174) & x(292) & x(293) & x(318) & x(321) & x(322) & x(327) & x(341) & x(342) & x(366) & x(369) & x(418) & x(426) & x(431) & x(459) & x(460) & x(472) & x(473) & x(475) & x(499) & x(507) & x(527) & x(584) & x(619) & x(697);
    y(161) <= not(p161_out);
    p161 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111001101000001000011111111111111",
            TABLE => "0000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101101110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 3,
            B => 49,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p161_in,
            y(0) => p161_out,
            y(1 to 14 - 1) => dummy161
        );


    p162_in <= x(35) & x(46) & x(63) & x(68) & x(69) & x(70) & x(73) & x(74) & x(78) & x(95) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(108) & x(190) & x(191) & x(192) & x(218) & x(219) & x(220) & x(221) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(278) & x(304) & x(305) & x(306) & x(307) & x(321) & x(329) & x(330) & x(333) & x(349) & x(359) & x(387) & x(388) & x(390) & x(415) & x(501) & x(529) & x(721) & x(746) & x(747);
    y(162) <= not(p162_out);
    p162 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111111111111110000000000000000000011001110111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => 49,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p162_in,
            y(0) => p162_out,
            y(1 to 14 - 1) => dummy162
        );


    p163_in <= x(40) & x(44) & x(64) & x(65) & x(66) & x(68) & x(91) & x(93) & x(94) & x(95) & x(96) & x(97) & x(99) & x(192) & x(220) & x(221) & x(238) & x(247) & x(248) & x(249) & x(267) & x(275) & x(276) & x(277) & x(278) & x(304) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(333) & x(334) & x(343) & x(357) & x(358) & x(359) & x(360) & x(371) & x(372) & x(387) & x(388) & x(396) & x(398) & x(399) & x(440) & x(445) & x(473) & x(501) & x(513) & x(514) & x(736) & x(740) & x(741) & x(742) & x(745) & x(746) & x(747);
    y(163) <= not(p163_out);
    p163 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111111110001000100000001111000111100110000111111111111",
            TABLE => "00000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100110110010001000000010000000000000111110111011001010110010001000001011001000100100001001000100110111011011101100101011001000100100100101100110100101101001100101100110100110010110100101100110100111101000111111101000000011101000100000001110100000000000100000001110100001111110100000011110100010000001111010000001011110000001011010011001011010010110011010011001011001101001011010011001011011110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100101000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011000000000010000000100000011010100010000001101010011010100111111010010101101000010010000101101010001000010110101001101010010111101100101100110100101101001100101100110100110010110100101100110100111010100010000000100000000000000111111011101010011010100010000001101010001000010010000100010101110111101110101001101010001000010100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000001000101110001011101111111100000010001011100010111011111100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 3,
            B => 71,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p163_in,
            y(0) => p163_out,
            y(1 to 15 - 1) => dummy163
        );


    p164_in <= x(35) & x(40) & x(46) & x(50) & x(64) & x(78) & x(91) & x(107) & x(108) & x(185) & x(186) & x(192) & x(210) & x(211) & x(212) & x(220) & x(239) & x(248) & x(249) & x(266) & x(267) & x(276) & x(277) & x(290) & x(292) & x(305) & x(306) & x(322) & x(328) & x(329) & x(330) & x(331) & x(332) & x(334) & x(350) & x(357) & x(358) & x(359) & x(360) & x(387) & x(388) & x(411) & x(415) & x(416) & x(438) & x(439) & x(446) & x(453) & x(566) & x(598) & x(719) & x(720) & x(746) & x(747);
    y(164) <= not(p164_out);
    p164 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000000001000101100111111000000100000001001110000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 2,
            B => -56,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p164_in,
            y(0) => p164_out,
            y(1 to 13 - 1) => dummy164
        );


    p165_in <= x(210) & x(220) & x(248) & x(275) & x(276) & x(277) & x(278) & x(284) & x(303) & x(304) & x(305) & x(306) & x(320) & x(333) & x(334) & x(361) & x(426) & x(427) & x(453) & x(454) & x(455) & x(584) & x(612) & x(668) & x(721) & x(732) & x(733);
    y(165) <= not(p165_out);
    p165 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011111111111111100000000000",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 3,
            B => 50,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p165_in,
            y(0) => p165_out,
            y(1 to 13 - 1) => dummy165
        );


    p166_in <= x(136) & x(165) & x(192) & x(193) & x(220) & x(221) & x(248) & x(249) & x(250) & x(274) & x(275) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(321) & x(322) & x(328) & x(329) & x(332) & x(333) & x(334) & x(348) & x(367) & x(455) & x(456) & x(479) & x(484) & x(485) & x(486) & x(487) & x(515) & x(685) & x(686) & x(746);
    y(166) <= not(p166_out);
    p166 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000000000110000011011111001",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 2,
            B => -83,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p166_in,
            y(0) => p166_out,
            y(1 to 13 - 1) => dummy166
        );


    p167_in <= x(145) & x(165) & x(172) & x(199) & x(200) & x(201) & x(220) & x(228) & x(248) & x(256) & x(275) & x(276) & x(277) & x(283) & x(289) & x(295) & x(303) & x(304) & x(305) & x(306) & x(310) & x(311) & x(323) & x(333) & x(334) & x(338) & x(339) & x(366) & x(368) & x(390) & x(402) & x(403) & x(418) & x(422) & x(430) & x(490) & x(500) & x(528) & x(535) & x(582) & x(667) & x(676) & x(677) & x(705) & x(708) & x(717) & x(724);
    y(167) <= not(p167_out);
    p167 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01000010101110101111000110000111101011011000011",
            TABLE => "11101000100000001111111011101000100000000000000011101000100000001110100010000001011111101110100010000001000101111110100010000001011010011001011010010110011010011001011001101001011010011001011000010000011100010000000000010000011100011111011100010000011100010001100001110001100011100001100001110001111001110001100001110001100101100110100101101001100101100110100110010110100101100110100100010000011100010000000000010000011100011111011100010000011100010001100001110001100011100001100001110001111001110001100001110001100101100110100101101001100101100110100110010110100101100110100101000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011011010100010000000100000000000000111111011101010011010100010000001101010001000010010000100010101110111101110101001101010001000010100101100110100101101001100101100110100110010110100101100110100100000000001000000010000010110010001000001011001010110010111110110100110100100100001001001011001000100100101100101011001011011011100101100110100101101001100101100110100110010110100101100110100100000010000000000010101100000010001010110000001010111111001010110100001011010100001010110100001000101011010000101011110100101011100101100110100101101001100101100110100110010110100101100110100111110111011100010111000100010000111001110111000101110001000110001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p167_in,
            y(0) => p167_out,
            y(1 to 14 - 1) => dummy167
        );


    p168_in <= x(162) & x(163) & x(192) & x(221) & x(222) & x(249) & x(277) & x(305) & x(311) & x(329) & x(330) & x(331) & x(332) & x(339) & x(357) & x(358) & x(359) & x(360) & x(386) & x(387) & x(388) & x(422) & x(427) & x(429) & x(430) & x(454) & x(455) & x(456) & x(457) & x(458) & x(483) & x(484) & x(485) & x(486) & x(487) & x(507) & x(515) & x(535) & x(659) & x(676) & x(681) & x(683) & x(684) & x(685) & x(686) & x(687) & x(708) & x(709) & x(710) & x(712) & x(769);
    y(168) <= not(p168_out);
    p168 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000000111101111111011111111111110100000000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 2,
            B => -35,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p168_in,
            y(0) => p168_out,
            y(1 to 13 - 1) => dummy168
        );


    p169_in <= x(67) & x(70) & x(71) & x(72) & x(73) & x(90) & x(91) & x(92) & x(93) & x(94) & x(97) & x(99) & x(118) & x(228) & x(248) & x(256) & x(276) & x(277) & x(283) & x(284) & x(285) & x(301) & x(304) & x(305) & x(310) & x(311) & x(312) & x(328) & x(339) & x(361) & x(366) & x(451) & x(479) & x(507) & x(535) & x(563) & x(619) & x(638) & x(639) & x(679) & x(694) & x(695) & x(732) & x(762);
    y(169) <= not(p169_out);
    p169 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000101100001100000000000001101110",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => -296,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p169_in,
            y(0) => p169_out,
            y(1 to 15 - 1) => dummy169
        );


    p170_in <= x(183) & x(222) & x(277) & x(302) & x(303) & x(305) & x(329) & x(330) & x(331) & x(332) & x(341) & x(342) & x(355) & x(357) & x(358) & x(359) & x(360) & x(387) & x(455) & x(473) & x(483) & x(501) & x(502) & x(528) & x(529) & x(556) & x(592) & x(620) & x(648) & x(649) & x(717) & x(719) & x(720) & x(746);
    y(170) <= not(p170_out);
    p170 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001101111111111111010000000001111",
            TABLE => "0010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 3,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p170_in,
            y(0) => p170_out,
            y(1 to 14 - 1) => dummy170
        );


    p171_in <= x(65) & x(78) & x(79) & x(80) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(102) & x(104) & x(108) & x(118) & x(148) & x(176) & x(186) & x(187) & x(200) & x(205) & x(228) & x(231) & x(248) & x(256) & x(257) & x(276) & x(277) & x(285) & x(286) & x(287) & x(304) & x(305) & x(310) & x(311) & x(312) & x(313) & x(328) & x(329) & x(330) & x(338) & x(339) & x(350) & x(356) & x(357) & x(359) & x(360) & x(366) & x(387) & x(417) & x(418) & x(445) & x(473) & x(501) & x(547) & x(548) & x(576) & x(604) & x(605) & x(619) & x(695) & x(697) & x(723);
    y(171) <= not(p171_out);
    p171 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000000000000001100001001100011000000000100000000000000000101",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001010011010110100111111111",
            SHIFT => 2,
            B => -162,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p171_in,
            y(0) => p171_out,
            y(1 to 14 - 1) => dummy171
        );


    p172_in <= x(97) & x(161) & x(190) & x(218) & x(353) & x(381) & x(408) & x(409) & x(416) & x(418) & x(437) & x(528) & x(542) & x(554) & x(557) & x(570) & x(571) & x(581) & x(586) & x(607) & x(609) & x(634) & x(635) & x(636) & x(637) & x(638) & x(697) & x(707) & x(711) & x(713) & x(714) & x(715) & x(719);
    y(172) <= not(p172_out);
    p172 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000011110010000000000000000111111",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => 2,
            B => -63,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p172_in,
            y(0) => p172_out,
            y(1 to 13 - 1) => dummy172
        );


    p173_in <= x(66) & x(68) & x(236) & x(247) & x(276) & x(277) & x(303) & x(304) & x(305) & x(306) & x(310) & x(332) & x(333) & x(338) & x(339) & x(366) & x(405) & x(432) & x(433) & x(450) & x(461) & x(611) & x(647) & x(720);
    y(173) <= not(p173_out);
    p173 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110011111101100011111011",
            TABLE => "000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => 47,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p173_in,
            y(0) => p173_out,
            y(1 to 13 - 1) => dummy173
        );


    p174_in <= x(40) & x(162) & x(198) & x(209) & x(228) & x(237) & x(263) & x(264) & x(299) & x(305) & x(328) & x(329) & x(330) & x(331) & x(332) & x(358) & x(359) & x(360) & x(361) & x(387) & x(388) & x(418) & x(443) & x(473) & x(501) & x(514) & x(529) & x(536) & x(584) & x(611) & x(638) & x(666) & x(696) & x(713) & x(743);
    y(174) <= not(p174_out);
    p174 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110111010000000000010110111111111",
            TABLE => "00000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100100001000000000001000111000001000100011100000100011101111100011100001100001110001100011100001100010001110000110001110011110001110011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111011111010011010100110100000100010011010000010000000100000000001101101101001101010011010010010001001101001001000010010010110010100101100110100101101001100101100110100110010110100101100110100100000001000101110000000000000001000101110111111100000001000101111000000100010111111010001000000100010111011111101000000100010111011010011001011010010110011010011001011001101001011010011001011000000001000101110001011101111111100000010001011100010111011111100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 3,
            B => 21,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p174_in,
            y(0) => p174_out,
            y(1 to 14 - 1) => dummy174
        );


    p175_in <= x(66) & x(71) & x(72) & x(73) & x(182) & x(192) & x(220) & x(228) & x(248) & x(249) & x(256) & x(276) & x(277) & x(297) & x(300) & x(304) & x(305) & x(306) & x(311) & x(328) & x(329) & x(330) & x(331) & x(332) & x(357) & x(358) & x(359) & x(360) & x(361) & x(387) & x(388) & x(389) & x(439) & x(446) & x(464) & x(492) & x(541) & x(543) & x(569) & x(571) & x(611);
    y(175) <= not(p175_out);
    p175 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000001001001100011111111111111111100000",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100110110010001000001111101110110010001000000000000010110010001000001011001000100100110110111011001000100100010011011011001000100100100101100110100101101001100101100110100110010110100101100110100110000000111010001110100011111110000000001000000010000000111010001000000111101000111010000111111000010111100000011000000111101000100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p175_in,
            y(0) => p175_out,
            y(1 to 14 - 1) => dummy175
        );


    p176_in <= x(116) & x(192) & x(220) & x(248) & x(249) & x(276) & x(277) & x(310) & x(338) & x(339) & x(342) & x(343) & x(347) & x(348) & x(349) & x(350) & x(362) & x(366) & x(370) & x(375) & x(376) & x(377) & x(389) & x(390) & x(391) & x(404) & x(418) & x(446) & x(474) & x(502) & x(529) & x(531) & x(557) & x(697) & x(741) & x(742) & x(745) & x(746) & x(774);
    y(176) <= not(p176_out);
    p176 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000011100000011000011101111111111111",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 3,
            B => 61,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p176_in,
            y(0) => p176_out,
            y(1 to 14 - 1) => dummy176
        );


    p177_in <= x(40) & x(49) & x(50) & x(69) & x(98) & x(99) & x(108) & x(211) & x(228) & x(255) & x(256) & x(310) & x(311) & x(331) & x(334) & x(338) & x(339) & x(359) & x(360) & x(366) & x(387) & x(388) & x(415) & x(416) & x(443) & x(444) & x(460) & x(469) & x(488) & x(667) & x(676) & x(677) & x(678) & x(690) & x(691) & x(692) & x(693) & x(694) & x(695) & x(704) & x(708) & x(720) & x(764);
    y(177) <= not(p177_out);
    p177 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111111011111101111111111101001110000001101",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101101011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => 172,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p177_in,
            y(0) => p177_out,
            y(1 to 14 - 1) => dummy177
        );


    p178_in <= x(40) & x(44) & x(95) & x(96) & x(98) & x(100) & x(171) & x(176) & x(241) & x(247) & x(297) & x(298) & x(304) & x(309) & x(338) & x(350) & x(357) & x(366) & x(378) & x(415) & x(418) & x(434) & x(444) & x(446) & x(462) & x(473) & x(495) & x(501) & x(529) & x(544) & x(557) & x(571) & x(691) & x(692) & x(705);
    y(178) <= not(p178_out);
    p178 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000011010010010000000110",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100110111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100110001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100111101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011010111111001010110010101100000010101111010010101100101011010000101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -177,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p178_in,
            y(0) => p178_out,
            y(1 to 14 - 1) => dummy178
        );


    p179_in <= x(65) & x(66) & x(90) & x(129) & x(130) & x(157) & x(158) & x(192) & x(199) & x(218) & x(220) & x(221) & x(228) & x(247) & x(248) & x(249) & x(275) & x(276) & x(277) & x(304) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(358) & x(359) & x(360) & x(376) & x(388) & x(399) & x(404) & x(418) & x(428) & x(437) & x(470) & x(473) & x(498) & x(508) & x(509) & x(510) & x(514) & x(525) & x(526) & x(528) & x(536) & x(538) & x(539) & x(548) & x(549) & x(550) & x(552) & x(553) & x(566) & x(567) & x(568) & x(569) & x(576) & x(578) & x(579) & x(584) & x(592) & x(595) & x(596) & x(597) & x(598) & x(599) & x(604) & x(605) & x(606) & x(607) & x(610) & x(611) & x(620) & x(632) & x(634) & x(649) & x(696) & x(697) & x(767);
    y(179) <= not(p179_out);
    p179 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000001000100000000011111110100001000000100000000000000000000000000000000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 1,
            B => -99,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p179_in,
            y(0) => p179_out,
            y(1 to 13 - 1) => dummy179
        );


    p180_in <= x(144) & x(145) & x(157) & x(165) & x(171) & x(191) & x(192) & x(199) & x(210) & x(218) & x(219) & x(220) & x(221) & x(231) & x(232) & x(234) & x(247) & x(248) & x(249) & x(260) & x(275) & x(276) & x(277) & x(278) & x(291) & x(292) & x(294) & x(295) & x(296) & x(305) & x(306) & x(307) & x(322) & x(323) & x(328) & x(329) & x(330) & x(331) & x(334) & x(350) & x(358) & x(359) & x(375) & x(378) & x(390) & x(403) & x(418) & x(446) & x(473) & x(500) & x(528) & x(583) & x(611) & x(626) & x(660) & x(694) & x(695) & x(705) & x(706) & x(708) & x(719) & x(720) & x(721) & x(733) & x(734) & x(735) & x(736) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(745) & x(746);
    y(180) <= not(p180_out);
    p180 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110010011000000000000000001110001111110111010000000000011111111111111111111",
            TABLE => "001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 2,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p180_in,
            y(0) => p180_out,
            y(1 to 14 - 1) => dummy180
        );


    p181_in <= x(64) & x(65) & x(66) & x(67) & x(68) & x(78) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(106) & x(122) & x(295) & x(305) & x(323) & x(331) & x(332) & x(357) & x(358) & x(359) & x(360) & x(361) & x(387) & x(388) & x(389) & x(396) & x(406) & x(445) & x(461) & x(512) & x(739);
    y(181) <= not(p181_out);
    p181 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000000000001110000000000110100",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010011000111000001000100011100001100010010110011010010000000000000000",
            SHIFT => 3,
            B => -154,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p181_in,
            y(0) => p181_out,
            y(1 to 14 - 1) => dummy181
        );


    p182_in <= x(95) & x(120) & x(125) & x(126) & x(127) & x(136) & x(159) & x(160) & x(186) & x(187) & x(188) & x(192) & x(220) & x(221) & x(228) & x(248) & x(249) & x(250) & x(256) & x(268) & x(269) & x(276) & x(277) & x(278) & x(297) & x(298) & x(299) & x(300) & x(304) & x(305) & x(306) & x(311) & x(326) & x(331) & x(333) & x(334) & x(338) & x(350) & x(359) & x(360) & x(366) & x(385) & x(387) & x(388) & x(406) & x(433) & x(501) & x(695) & x(719) & x(723);
    y(182) <= not(p182_out);
    p182 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000111111111011100011100001110001101000100110111",
            TABLE => "111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 2,
            B => 42,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p182_in,
            y(0) => p182_out,
            y(1 to 13 - 1) => dummy182
        );


    p183_in <= x(220) & x(247) & x(248) & x(249) & x(275) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(333) & x(334) & x(362) & x(718) & x(745);
    y(183) <= not(p183_out);
    p183 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000000000",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -250,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p183_in,
            y(0) => p183_out,
            y(1 to 14 - 1) => dummy183
        );


    p184_in <= x(64) & x(66) & x(91) & x(92) & x(93) & x(95) & x(189) & x(206) & x(207) & x(213) & x(214) & x(215) & x(216) & x(235) & x(241) & x(242) & x(243) & x(305) & x(309) & x(310) & x(334) & x(338) & x(354) & x(359) & x(366) & x(387) & x(388) & x(415) & x(416) & x(418) & x(433) & x(434) & x(435) & x(444) & x(461) & x(462) & x(482) & x(489) & x(507) & x(599) & x(691) & x(704) & x(705) & x(707) & x(708) & x(747);
    y(184) <= not(p184_out);
    p184 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000000000000010010100000001110110110100000",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101101011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101101110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 2,
            B => -67,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p184_in,
            y(0) => p184_out,
            y(1 to 13 - 1) => dummy184
        );


    p185_in <= x(44) & x(104) & x(105) & x(106) & x(134) & x(135) & x(159) & x(160) & x(161) & x(162) & x(163) & x(164) & x(191) & x(192) & x(198) & x(221) & x(222) & x(249) & x(265) & x(269) & x(277) & x(299) & x(305) & x(309) & x(330) & x(331) & x(332) & x(338) & x(361) & x(362) & x(366) & x(374) & x(377) & x(378) & x(389) & x(390) & x(391) & x(400) & x(401) & x(406) & x(413) & x(414) & x(418) & x(446) & x(474) & x(475) & x(485) & x(500) & x(555) & x(583) & x(676) & x(694) & x(745) & x(746) & x(747) & x(774);
    y(185) <= not(p185_out);
    p185 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01111111111111011100101000000001110001111100000000110000",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 3,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p185_in,
            y(0) => p185_out,
            y(1 to 14 - 1) => dummy185
        );


    p186_in <= x(64) & x(66) & x(68) & x(91) & x(93) & x(108) & x(192) & x(214) & x(276) & x(277) & x(305) & x(328) & x(329) & x(330) & x(331) & x(332) & x(334) & x(356) & x(357) & x(358) & x(359) & x(360) & x(386) & x(387) & x(388) & x(417) & x(535) & x(546) & x(547) & x(574) & x(575) & x(602) & x(720) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(746);
    y(186) <= not(p186_out);
    p186 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111110000011111011111111101111111111111",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 2,
            B => 96,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p186_in,
            y(0) => p186_out,
            y(1 to 13 - 1) => dummy186
        );


    p187_in <= x(98) & x(276) & x(277) & x(293) & x(303) & x(304) & x(305) & x(306) & x(331) & x(332) & x(333) & x(334) & x(345) & x(387) & x(414) & x(415) & x(416) & x(442) & x(443) & x(444) & x(469) & x(471);
    y(187) <= not(p187_out);
    p187 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110111111111111111111",
            TABLE => "0000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 3,
            B => 135,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p187_in,
            y(0) => p187_out,
            y(1 to 13 - 1) => dummy187
        );


    p188_in <= x(66) & x(136) & x(249) & x(276) & x(277) & x(304) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(333) & x(334) & x(357) & x(358) & x(359) & x(360) & x(403) & x(425) & x(453) & x(454) & x(455) & x(461) & x(475) & x(481) & x(482) & x(483) & x(509) & x(510) & x(511) & x(512) & x(538) & x(539) & x(547) & x(566) & x(567) & x(574) & x(575) & x(602) & x(653) & x(675) & x(677) & x(678) & x(679) & x(680) & x(685) & x(686) & x(709) & x(746);
    y(188) <= not(p188_out);
    p188 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000111100111111111011111111111111110000000001",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 2,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p188_in,
            y(0) => p188_out,
            y(1 to 13 - 1) => dummy188
        );


    p189_in <= x(41) & x(183) & x(201) & x(203) & x(205) & x(231) & x(310) & x(311) & x(312) & x(339) & x(344) & x(345) & x(366) & x(370) & x(378) & x(387) & x(388) & x(397) & x(399) & x(405) & x(414) & x(415) & x(416) & x(422) & x(433) & x(441) & x(442) & x(443) & x(450) & x(466) & x(493) & x(535) & x(676) & x(692) & x(695) & x(704) & x(720);
    y(189) <= not(p189_out);
    p189 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1011111111111101111011110111111110010",
            TABLE => "0000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 2,
            B => 95,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p189_in,
            y(0) => p189_out,
            y(1 to 13 - 1) => dummy189
        );


    p190_in <= x(228) & x(256) & x(311) & x(341) & x(342) & x(343) & x(349) & x(358) & x(359) & x(360) & x(369) & x(370) & x(386) & x(387) & x(388) & x(390) & x(418) & x(446) & x(473) & x(474) & x(501) & x(502) & x(529);
    y(190) <= not(p190_out);
    p190 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11100000000000011111111",
            TABLE => "00000000100000001000000011101000100000001110100011101000111111100001011110000001100000011110100010000001111010001110100001111110011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100101111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011000000001000101110001011101111111100000010001011100010111011111100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 3,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p190_in,
            y(0) => p190_out,
            y(1 to 13 - 1) => dummy190
        );


    p191_in <= x(35) & x(65) & x(66) & x(68) & x(71) & x(91) & x(93) & x(100) & x(108) & x(210) & x(212) & x(213) & x(248) & x(276) & x(277) & x(285) & x(304) & x(305) & x(310) & x(312) & x(333) & x(334) & x(338) & x(339) & x(359) & x(360) & x(366) & x(369) & x(387) & x(388) & x(389) & x(462) & x(473) & x(490) & x(516) & x(517) & x(518) & x(519) & x(543) & x(544) & x(545) & x(546) & x(547) & x(572) & x(573) & x(659) & x(675) & x(694) & x(695) & x(697) & x(705) & x(720) & x(732) & x(751);
    y(191) <= not(p191_out);
    p191 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111000000100110011111011111111111111111100010000",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 2,
            B => 31,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p191_in,
            y(0) => p191_out,
            y(1 to 13 - 1) => dummy191
        );


    p192_in <= x(66) & x(70) & x(76) & x(105) & x(247) & x(248) & x(249) & x(276) & x(277) & x(305) & x(331) & x(359) & x(360) & x(388) & x(389) & x(391) & x(396) & x(473);
    y(192) <= not(p192_out);
    p192 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000011111100000010",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -82,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p192_in,
            y(0) => p192_out,
            y(1 to 14 - 1) => dummy192
        );


    p193_in <= x(40) & x(44) & x(109) & x(218) & x(245) & x(274) & x(277) & x(304) & x(305) & x(306) & x(375) & x(414) & x(415) & x(416) & x(434) & x(443) & x(444) & x(446) & x(470) & x(471) & x(472) & x(479) & x(480) & x(486) & x(487) & x(488) & x(489) & x(498) & x(508) & x(509) & x(515) & x(525) & x(526) & x(527) & x(537) & x(564) & x(569) & x(570) & x(571) & x(592) & x(640) & x(647) & x(720);
    y(193) <= not(p193_out);
    p193 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000000000010000000011110001000000000101",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101101111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101101110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 2,
            B => -110,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p193_in,
            y(0) => p193_out,
            y(1 to 13 - 1) => dummy193
        );


    p194_in <= x(248) & x(255) & x(275) & x(276) & x(277) & x(305) & x(306) & x(315) & x(316) & x(350) & x(359) & x(390) & x(391) & x(539) & x(582) & x(583) & x(584) & x(608) & x(610) & x(611) & x(636) & x(638) & x(665) & x(666) & x(697);
    y(194) <= not(p194_out);
    p194 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100000001100000000000000",
            TABLE => "1110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101101011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -203,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p194_in,
            y(0) => p194_out,
            y(1 to 14 - 1) => dummy194
        );


    p195_in <= x(116) & x(247) & x(248) & x(249) & x(276) & x(277) & x(304) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(357) & x(358) & x(359) & x(360) & x(366) & x(508) & x(528) & x(556) & x(557) & x(568) & x(570) & x(611) & x(695) & x(697);
    y(195) <= not(p195_out);
    p195 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011111111000000001111111101",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001010011010110100111111111",
            SHIFT => 3,
            B => 82,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p195_in,
            y(0) => p195_out,
            y(1 to 13 - 1) => dummy195
        );


    p196_in <= x(190) & x(192) & x(193) & x(219) & x(221) & x(249) & x(250) & x(276) & x(277) & x(305) & x(306) & x(318) & x(319) & x(320) & x(325) & x(333) & x(345) & x(351) & x(352) & x(353) & x(366) & x(380) & x(418) & x(422) & x(424) & x(425) & x(428) & x(446) & x(474) & x(475) & x(502) & x(507) & x(528) & x(546) & x(547) & x(557) & x(583) & x(611) & x(636) & x(637) & x(669) & x(679) & x(697) & x(705) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(713) & x(715) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(745) & x(749) & x(750);
    y(196) <= not(p196_out);
    p196 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011011111111111111111101000000010000000001011111111111111111111",
            TABLE => "000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 3,
            B => 91,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p196_in,
            y(0) => p196_out,
            y(1 to 15 - 1) => dummy196
        );


    p197_in <= x(66) & x(78) & x(91) & x(93) & x(101) & x(102) & x(103) & x(104) & x(106) & x(107) & x(108) & x(186) & x(187) & x(188) & x(189) & x(190) & x(192) & x(213) & x(214) & x(215) & x(216) & x(218) & x(228) & x(240) & x(242) & x(248) & x(256) & x(276) & x(277) & x(305) & x(306) & x(327) & x(334) & x(338) & x(359) & x(360) & x(366) & x(387) & x(388) & x(396) & x(575) & x(694) & x(695);
    y(197) <= not(p197_out);
    p197 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111111111100000000000100010000101111110100",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101101110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010010000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 2,
            B => 20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p197_in,
            y(0) => p197_out,
            y(1 to 13 - 1) => dummy197
        );


    p198_in <= x(95) & x(161) & x(162) & x(192) & x(220) & x(221) & x(247) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(317) & x(321) & x(322) & x(328) & x(333) & x(366) & x(458) & x(705);
    y(198) <= not(p198_out);
    p198 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01111111111111111111101100",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 3,
            B => 156,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p198_in,
            y(0) => p198_out,
            y(1 to 13 - 1) => dummy198
        );


    p199_in <= x(118) & x(121) & x(122) & x(123) & x(124) & x(125) & x(126) & x(127) & x(147) & x(286) & x(305) & x(311) & x(319) & x(333) & x(345) & x(347) & x(358) & x(359) & x(362) & x(373) & x(374) & x(375) & x(387) & x(388) & x(389) & x(390) & x(391) & x(418) & x(446) & x(451) & x(461) & x(474) & x(475) & x(488) & x(502) & x(531) & x(557) & x(558) & x(583) & x(584) & x(611) & x(619) & x(629) & x(638) & x(649) & x(744) & x(772);
    y(199) <= not(p199_out);
    p199 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000000000010111101111100000000000000000010000",
            TABLE => "11111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100000001000101110000000000000001000101110111111100000001000101111000000100010111111010001000000100010111011111101000000100010111011010011001011010010110011010011001011001101001011010011001011000000001000101110001011101111111000000000000000100000001000101111000000100010111000101110111111011101000100000011000000100010111011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111101000100000001111111011101000111010001000000101111110111010000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 2,
            B => -138,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p199_in,
            y(0) => p199_out,
            y(1 to 13 - 1) => dummy199
        );


    p200_in <= x(93) & x(95) & x(96) & x(108) & x(249) & x(276) & x(277) & x(305) & x(313) & x(323) & x(331) & x(333) & x(334) & x(340) & x(341) & x(342) & x(358) & x(359) & x(360) & x(368) & x(369) & x(374) & x(387) & x(388) & x(389) & x(396) & x(399) & x(400) & x(401) & x(403) & x(415) & x(416) & x(429) & x(442) & x(443) & x(444) & x(445) & x(470) & x(471) & x(473) & x(498) & x(501) & x(517) & x(529) & x(717) & x(719) & x(720) & x(721);
    y(200) <= not(p200_out);
    p200 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111100000010000011100111101111111111111111010000",
            TABLE => "000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 2,
            B => 21,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p200_in,
            y(0) => p200_out,
            y(1 to 13 - 1) => dummy200
        );


    p201_in <= x(62) & x(63) & x(65) & x(66) & x(72) & x(73) & x(90) & x(91) & x(93) & x(102) & x(105) & x(182) & x(249) & x(250) & x(277) & x(305) & x(306) & x(331) & x(359) & x(360) & x(387) & x(388) & x(396) & x(397) & x(415) & x(416) & x(424) & x(442) & x(443) & x(529) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(737) & x(738) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(748) & x(750);
    y(201) <= not(p201_out);
    p201 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111111111110000000000001111111111111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => 205,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p201_in,
            y(0) => p201_out,
            y(1 to 14 - 1) => dummy201
        );


    p202_in <= x(66) & x(106) & x(192) & x(220) & x(221) & x(247) & x(248) & x(249) & x(276) & x(277) & x(302) & x(305) & x(328) & x(329) & x(330) & x(331) & x(418) & x(424) & x(425) & x(446) & x(452) & x(453) & x(474) & x(502);
    y(202) <= not(p202_out);
    p202 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000000010111111111111",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => 23,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p202_in,
            y(0) => p202_out,
            y(1 to 13 - 1) => dummy202
        );


    p203_in <= x(35) & x(62) & x(63) & x(64) & x(66) & x(68) & x(69) & x(90) & x(91) & x(92) & x(95) & x(101) & x(102) & x(103) & x(104) & x(106) & x(108) & x(220) & x(230) & x(231) & x(242) & x(247) & x(248) & x(269) & x(271) & x(276) & x(284) & x(298) & x(299) & x(307) & x(309) & x(310) & x(313) & x(314) & x(338) & x(366) & x(374) & x(401) & x(402) & x(573) & x(574) & x(659) & x(660) & x(661) & x(668) & x(694) & x(695) & x(720) & x(732) & x(733);
    y(203) <= not(p203_out);
    p203 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111111111111000000000000000000011111000111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 2,
            B => 42,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p203_in,
            y(0) => p203_out,
            y(1 to 13 - 1) => dummy203
        );


    p204_in <= x(62) & x(63) & x(64) & x(65) & x(66) & x(135) & x(228) & x(229) & x(276) & x(277) & x(300) & x(302) & x(304) & x(305) & x(306) & x(330) & x(331) & x(332) & x(359) & x(360) & x(361) & x(406) & x(407) & x(455) & x(501) & x(528) & x(544) & x(611) & x(666) & x(718) & x(724);
    y(204) <= not(p204_out);
    p204 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000001100110001111110010000000",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => -68,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p204_in,
            y(0) => p204_out,
            y(1 to 14 - 1) => dummy204
        );


    p205_in <= x(95) & x(96) & x(98) & x(171) & x(192) & x(220) & x(248) & x(266) & x(267) & x(277) & x(294) & x(295) & x(296) & x(309) & x(310) & x(311) & x(338) & x(339) & x(358) & x(366) & x(384) & x(385) & x(391) & x(418) & x(474) & x(475) & x(501) & x(502) & x(529) & x(557) & x(667) & x(676) & x(692) & x(695) & x(705) & x(706) & x(708) & x(742) & x(745) & x(746) & x(747) & x(750);
    y(205) <= not(p205_out);
    p205 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000011100100000000101100000000101100000000",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => -130,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p205_in,
            y(0) => p205_out,
            y(1 to 14 - 1) => dummy205
        );


    p206_in <= x(136) & x(192) & x(198) & x(221) & x(236) & x(248) & x(249) & x(268) & x(269) & x(276) & x(277) & x(297) & x(298) & x(299) & x(304) & x(305) & x(306) & x(309) & x(310) & x(333) & x(334) & x(338) & x(349) & x(350) & x(366) & x(418) & x(435) & x(446) & x(474) & x(485) & x(501) & x(507) & x(583) & x(675) & x(694) & x(695) & x(720) & x(723) & x(774);
    y(206) <= not(p206_out);
    p206 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001010011001110001100100110111101000001",
            TABLE => "101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001110101001001011011111111",
            SHIFT => 3,
            B => -41,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p206_in,
            y(0) => p206_out,
            y(1 to 14 - 1) => dummy206
        );


    p207_in <= x(66) & x(183) & x(192) & x(220) & x(221) & x(248) & x(249) & x(276) & x(277) & x(304) & x(305) & x(306) & x(320) & x(321) & x(329) & x(330) & x(348) & x(357) & x(358) & x(474) & x(486) & x(513) & x(514) & x(515) & x(742);
    y(207) <= not(p207_out);
    p207 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100000000000011011111111",
            TABLE => "1110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010100110111011111000001000100110100000100010011010000000000000100010011011101101100100100010011010010010001001101101100100010010001101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => -30,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p207_in,
            y(0) => p207_out,
            y(1 to 13 - 1) => dummy207
        );


    p208_in <= x(35) & x(62) & x(64) & x(65) & x(67) & x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(76) & x(79) & x(80) & x(90) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(97) & x(99) & x(100) & x(101) & x(102) & x(103) & x(104) & x(105) & x(108) & x(118) & x(122) & x(192) & x(198) & x(228) & x(231) & x(248) & x(249) & x(256) & x(266) & x(276) & x(277) & x(304) & x(305) & x(310) & x(318) & x(328) & x(329) & x(330) & x(331) & x(332) & x(334) & x(338) & x(339) & x(358) & x(359) & x(360) & x(361) & x(366) & x(375) & x(387) & x(388) & x(389) & x(396) & x(397) & x(417) & x(418) & x(432) & x(473) & x(474) & x(707) & x(708) & x(735) & x(736) & x(739) & x(741) & x(742) & x(744) & x(745) & x(746) & x(747) & x(764) & x(769) & x(770);
    y(208) <= not(p208_out);
    p208 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111111111111111111111111111110111001100001011111011111110111001101111111111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 3,
            B => 362,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p208_in,
            y(0) => p208_out,
            y(1 to 15 - 1) => dummy208
        );


    p209_in <= x(69) & x(70) & x(106) & x(171) & x(209) & x(237) & x(247) & x(248) & x(249) & x(269) & x(276) & x(277) & x(304) & x(305) & x(306) & x(307) & x(309) & x(310) & x(329) & x(330) & x(338) & x(357) & x(358) & x(359) & x(360) & x(362) & x(366) & x(379) & x(384) & x(385) & x(387) & x(389) & x(390) & x(391) & x(418) & x(434) & x(446) & x(462) & x(473) & x(474) & x(500) & x(501) & x(502) & x(528) & x(557);
    y(209) <= not(p209_out);
    p209 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111000000000000000110111100111100001010000000",
            TABLE => "000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 3,
            B => -115,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p209_in,
            y(0) => p209_out,
            y(1 to 14 - 1) => dummy209
        );


    p210_in <= x(95) & x(98) & x(267) & x(277) & x(294) & x(295) & x(305) & x(321) & x(322) & x(390) & x(611) & x(665) & x(745) & x(746) & x(747);
    y(210) <= not(p210_out);
    p210 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111011011000111",
            TABLE => "000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 3,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p210_in,
            y(0) => p210_out,
            y(1 to 13 - 1) => dummy210
        );


    p211_in <= x(106) & x(236) & x(237) & x(241) & x(255) & x(266) & x(309) & x(310) & x(333) & x(338) & x(339) & x(357) & x(358) & x(366) & x(374) & x(375) & x(398) & x(399) & x(400) & x(401) & x(403) & x(426) & x(427) & x(428) & x(454) & x(456) & x(458) & x(484) & x(501) & x(611) & x(637) & x(664) & x(665) & x(666) & x(669) & x(677) & x(678) & x(685) & x(693) & x(706) & x(707) & x(708) & x(709) & x(711) & x(712) & x(714) & x(715) & x(718) & x(719) & x(724) & x(732) & x(739) & x(741) & x(743) & x(744) & x(745) & x(747) & x(748) & x(750) & x(764) & x(769) & x(774);
    y(211) <= not(p211_out);
    p211 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01111111111001000000000000000000000111011111111111011111111111",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 2,
            B => 55,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p211_in,
            y(0) => p211_out,
            y(1 to 14 - 1) => dummy211
        );


    p212_in <= x(63) & x(64) & x(65) & x(66) & x(67) & x(145) & x(159) & x(160) & x(174) & x(199) & x(201) & x(228) & x(256) & x(276) & x(277) & x(283) & x(296) & x(297) & x(299) & x(301) & x(302) & x(304) & x(305) & x(306) & x(310) & x(311) & x(330) & x(331) & x(338) & x(339) & x(359) & x(360) & x(361) & x(366) & x(378) & x(388) & x(405) & x(406) & x(422) & x(528) & x(582) & x(638) & x(666) & x(668) & x(679) & x(767);
    y(212) <= not(p212_out);
    p212 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111101100000110000001110000000000101101111101",
            TABLE => "0000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100000010001001101001001000100110110010110011010010000000000000000",
            SHIFT => 3,
            B => -30,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p212_in,
            y(0) => p212_out,
            y(1 to 14 - 1) => dummy212
        );


    p213_in <= x(93) & x(106) & x(108) & x(171) & x(176) & x(248) & x(250) & x(276) & x(277) & x(305) & x(306) & x(321) & x(333) & x(342) & x(438) & x(439) & x(462) & x(466) & x(490) & x(516) & x(705) & x(706) & x(707);
    y(213) <= not(p213_out);
    p213 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00011111111111110100111",
            TABLE => "01111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000001000000010001001101000001000100110101001101110111111011001000100100001001000100110100100100010011010100110111011011011010011001011010010110011010011001011001101001011010011001011001111111000101110001011100000001011111100001011100010111100000010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 3,
            B => 83,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p213_in,
            y(0) => p213_out,
            y(1 to 13 - 1) => dummy213
        );


    p214_in <= x(44) & x(65) & x(67) & x(144) & x(145) & x(171) & x(198) & x(306) & x(311) & x(334) & x(368) & x(369) & x(370) & x(371) & x(389) & x(390) & x(396) & x(397) & x(398) & x(418) & x(424) & x(425) & x(426) & x(442) & x(446) & x(473) & x(474) & x(500) & x(501) & x(528) & x(529) & x(676) & x(705) & x(717);
    y(214) <= not(p214_out);
    p214 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001110010111100111011110000000110",
            TABLE => "0111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101100001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010010000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 3,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p214_in,
            y(0) => p214_out,
            y(1 to 14 - 1) => dummy214
        );


    p215_in <= x(136) & x(185) & x(205) & x(206) & x(222) & x(232) & x(233) & x(240) & x(260) & x(261) & x(288) & x(289) & x(295) & x(311) & x(314) & x(315) & x(316) & x(319) & x(341) & x(342) & x(343) & x(358) & x(369) & x(418) & x(473) & x(501) & x(502) & x(529) & x(545) & x(582) & x(629) & x(657) & x(690) & x(705);
    y(215) <= not(p215_out);
    p215 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000100000001100000000011111100001",
            TABLE => "1111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101101010001000000110101000100001010010110011010010000000000000000",
            SHIFT => 2,
            B => -17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p215_in,
            y(0) => p215_out,
            y(1 to 13 - 1) => dummy215
        );


    p216_in <= x(68) & x(69) & x(70) & x(71) & x(72) & x(73) & x(74) & x(75) & x(91) & x(92) & x(93) & x(94) & x(95) & x(96) & x(102) & x(108) & x(171) & x(199) & x(228) & x(248) & x(276) & x(277) & x(305) & x(310) & x(328) & x(329) & x(330) & x(332) & x(338) & x(339) & x(366) & x(374) & x(396) & x(401) & x(402) & x(403) & x(609) & x(621) & x(623) & x(637) & x(638) & x(648) & x(649) & x(650) & x(651) & x(652) & x(665) & x(677) & x(678) & x(679) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(745) & x(774);
    y(216) <= not(p216_out);
    p216 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000000000000000111100000000111111001100000100000000000",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101101111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 3,
            B => -210,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p216_in,
            y(0) => p216_out,
            y(1 to 14 - 1) => dummy216
        );


    p217_in <= x(145) & x(156) & x(157) & x(180) & x(205) & x(206) & x(233) & x(244) & x(247) & x(248) & x(260) & x(276) & x(277) & x(305) & x(306) & x(314) & x(315) & x(329) & x(330) & x(351) & x(378) & x(406) & x(407) & x(434) & x(435) & x(461) & x(462) & x(473) & x(489) & x(490) & x(501) & x(516) & x(517) & x(540) & x(541) & x(609) & x(635) & x(657) & x(658) & x(659) & x(688);
    y(217) <= not(p217_out);
    p217 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000000000000000111111111111111100000000",
            TABLE => "11101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111101110101001101010001000000110101000100000001000000000000001011110111010100110101000100001011010100010000100100001000101011011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000100000001000000011101000100000001110100011101000111111100001011110000001100000011110100010000001111010001110100001111110011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 2,
            B => -24,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p217_in,
            y(0) => p217_out,
            y(1 to 13 - 1) => dummy217
        );


    p218_in <= x(95) & x(98) & x(99) & x(100) & x(101) & x(108) & x(118) & x(120) & x(136) & x(183) & x(184) & x(185) & x(211) & x(212) & x(213) & x(220) & x(248) & x(276) & x(277) & x(305) & x(306) & x(311) & x(333) & x(334) & x(360) & x(379) & x(387) & x(388) & x(399) & x(415) & x(416) & x(418) & x(424) & x(425) & x(426) & x(427) & x(454) & x(469) & x(501) & x(502) & x(529) & x(535) & x(557) & x(558) & x(564) & x(619) & x(676) & x(691) & x(692) & x(695) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(769) & x(772);
    y(218) <= not(p218_out);
    p218 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111110000000000000100101111111111111111111110000000000011",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 2,
            B => 65,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p218_in,
            y(0) => p218_out,
            y(1 to 14 - 1) => dummy218
        );


    p219_in <= x(117) & x(145) & x(171) & x(249) & x(277) & x(294) & x(305) & x(311) & x(321) & x(322) & x(323) & x(333) & x(339) & x(358) & x(359) & x(366) & x(387) & x(390) & x(391) & x(451) & x(479) & x(620) & x(621) & x(648) & x(649) & x(650) & x(651) & x(676) & x(677) & x(705) & x(706) & x(707) & x(708) & x(709) & x(736) & x(737) & x(744) & x(745) & x(746) & x(750) & x(772) & x(773);
    y(219) <= not(p219_out);
    p219 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111111100101111111111111111111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => 239,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p219_in,
            y(0) => p219_out,
            y(1 to 14 - 1) => dummy219
        );


    p220_in <= x(70) & x(71) & x(73) & x(74) & x(102) & x(131) & x(149) & x(173) & x(174) & x(177) & x(192) & x(193) & x(201) & x(204) & x(205) & x(206) & x(221) & x(233) & x(234) & x(243) & x(249) & x(270) & x(273) & x(274) & x(276) & x(277) & x(284) & x(301) & x(305) & x(306) & x(322) & x(330) & x(331) & x(334) & x(350) & x(358) & x(359) & x(360) & x(378) & x(387) & x(405) & x(406) & x(434) & x(480) & x(486) & x(492) & x(507) & x(508) & x(509) & x(514) & x(515) & x(527) & x(537) & x(543) & x(544) & x(553) & x(565) & x(572) & x(580) & x(584) & x(606) & x(607) & x(608) & x(611) & x(620) & x(634) & x(635) & x(636) & x(637) & x(662) & x(663) & x(664) & x(665) & x(685) & x(710);
    y(220) <= not(p220_out);
    p220 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000111111111111111111111111000100000000010111100110011011111111111111111",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 2,
            B => 62,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p220_in,
            y(0) => p220_out,
            y(1 to 14 - 1) => dummy220
        );


    p221_in <= x(74) & x(75) & x(192) & x(198) & x(208) & x(209) & x(210) & x(211) & x(212) & x(220) & x(221) & x(238) & x(248) & x(249) & x(250) & x(276) & x(277) & x(278) & x(305) & x(306) & x(328) & x(329) & x(333) & x(334) & x(338) & x(366) & x(418) & x(426) & x(453) & x(454) & x(474) & x(475) & x(501) & x(508) & x(584) & x(612) & x(640) & x(668) & x(697) & x(713) & x(714) & x(715) & x(741) & x(742) & x(743) & x(745) & x(746) & x(774);
    y(221) <= not(p221_out);
    p221 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111000000110111111110011000000000000000000000000",
            TABLE => "000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => -59,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p221_in,
            y(0) => p221_out,
            y(1 to 14 - 1) => dummy221
        );


    p222_in <= x(44) & x(98) & x(99) & x(100) & x(171) & x(192) & x(199) & x(202) & x(208) & x(227) & x(228) & x(236) & x(241) & x(242) & x(243) & x(248) & x(255) & x(256) & x(266) & x(267) & x(277) & x(283) & x(294) & x(295) & x(296) & x(309) & x(310) & x(311) & x(317) & x(334) & x(338) & x(339) & x(358) & x(366) & x(385) & x(418) & x(433) & x(529) & x(557) & x(613) & x(665) & x(667) & x(676) & x(677) & x(678) & x(691) & x(692) & x(695) & x(704) & x(705) & x(706) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(713) & x(736) & x(737) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(750) & x(764) & x(773) & x(774);
    y(222) <= not(p222_out);
    p222 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111110111111111011110111111100110101011100111000111111111111111111111111",
            TABLE => "000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 2,
            B => 200,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p222_in,
            y(0) => p222_out,
            y(1 to 14 - 1) => dummy222
        );


    p223_in <= x(44) & x(122) & x(133) & x(134) & x(135) & x(159) & x(162) & x(163) & x(188) & x(189) & x(190) & x(191) & x(192) & x(217) & x(219) & x(220) & x(238) & x(248) & x(249) & x(276) & x(277) & x(305) & x(320) & x(322) & x(330) & x(331) & x(332) & x(342) & x(343) & x(344) & x(348) & x(350) & x(357) & x(358) & x(360) & x(370) & x(389) & x(390) & x(391) & x(396) & x(418) & x(446) & x(473) & x(474) & x(475) & x(501) & x(502) & x(520) & x(529) & x(650) & x(653) & x(661) & x(666) & x(668) & x(678) & x(679) & x(680) & x(681) & x(697) & x(713) & x(714) & x(732) & x(733) & x(738);
    y(223) <= not(p223_out);
    p223 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0011111111111111011111110001111100010001000000000111001111000000",
            TABLE => "0001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101101110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010011110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 2,
            B => 21,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p223_in,
            y(0) => p223_out,
            y(1 to 14 - 1) => dummy223
        );


    p224_in <= x(66) & x(68) & x(70) & x(160) & x(161) & x(162) & x(183) & x(192) & x(221) & x(249) & x(276) & x(277) & x(287) & x(304) & x(305) & x(306) & x(310) & x(312) & x(314) & x(330) & x(331) & x(339) & x(358) & x(359) & x(366) & x(459) & x(484) & x(486) & x(513) & x(536) & x(592) & x(620) & x(648) & x(649) & x(653) & x(677) & x(769);
    y(224) <= not(p224_out);
    p224 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000001000000000000110110111100000000",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => -197,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p224_in,
            y(0) => p224_out,
            y(1 to 14 - 1) => dummy224
        );


    p225_in <= x(35) & x(46) & x(62) & x(63) & x(64) & x(66) & x(68) & x(78) & x(91) & x(106) & x(107) & x(108) & x(132) & x(133) & x(134) & x(135) & x(156) & x(161) & x(162) & x(163) & x(368) & x(390) & x(446) & x(485) & x(705) & x(721) & x(734) & x(738) & x(739) & x(740) & x(741) & x(742) & x(743) & x(746);
    y(225) <= not(p225_out);
    p225 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000000000000100001110000000000",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 4,
            B => -389,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p225_in,
            y(0) => p225_out,
            y(1 to 15 - 1) => dummy225
        );


    p226_in <= x(98) & x(123) & x(127) & x(128) & x(129) & x(151) & x(153) & x(155) & x(156) & x(157) & x(178) & x(179) & x(180) & x(181) & x(182) & x(227) & x(228) & x(248) & x(256) & x(276) & x(277) & x(305) & x(310) & x(312) & x(338) & x(339) & x(340) & x(358) & x(359) & x(360) & x(366) & x(375) & x(387) & x(388) & x(403) & x(430) & x(498) & x(516) & x(521) & x(523) & x(525) & x(538) & x(548) & x(549) & x(551) & x(566) & x(569) & x(580) & x(638);
    y(226) <= not(p226_out);
    p226 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111111111111110010111000000000100111011111111111",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010010000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101100000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 2,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p226_in,
            y(0) => p226_out,
            y(1 to 13 - 1) => dummy226
        );


    p227_in <= x(136) & x(192) & x(198) & x(221) & x(228) & x(236) & x(238) & x(248) & x(249) & x(256) & x(264) & x(265) & x(266) & x(276) & x(277) & x(294) & x(302) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(332) & x(338) & x(347) & x(348) & x(357) & x(358) & x(359) & x(360) & x(361) & x(366) & x(375) & x(376) & x(387) & x(388) & x(389) & x(391) & x(418) & x(454) & x(515) & x(546) & x(613) & x(675) & x(715) & x(716) & x(718) & x(720) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(774);
    y(227) <= not(p227_out);
    p227 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101000110000110011000000110000001100000000010000000000000",
            TABLE => "0000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101101000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101101110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010011011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 2,
            B => -95,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p227_in,
            y(0) => p227_out,
            y(1 to 14 - 1) => dummy227
        );


    p228_in <= x(95) & x(96) & x(98) & x(106) & x(122) & x(124) & x(150) & x(163) & x(171) & x(192) & x(220) & x(228) & x(248) & x(255) & x(270) & x(271) & x(277) & x(295) & x(296) & x(297) & x(298) & x(299) & x(300) & x(309) & x(310) & x(311) & x(316) & x(317) & x(325) & x(326) & x(338) & x(339) & x(366) & x(376) & x(377) & x(378) & x(535) & x(557) & x(665) & x(676) & x(690) & x(692) & x(704) & x(705) & x(708) & x(774);
    y(228) <= not(p228_out);
    p228 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110111010010111011111111100111110001101001111",
            TABLE => "0000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010010000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101100000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 2,
            B => 63,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p228_in,
            y(0) => p228_out,
            y(1 to 13 - 1) => dummy228
        );


    p229_in <= x(35) & x(41) & x(78) & x(269) & x(338) & x(350) & x(366) & x(379) & x(380) & x(390) & x(391) & x(418) & x(446) & x(480) & x(481) & x(482) & x(508) & x(509) & x(510) & x(528) & x(531) & x(536) & x(555) & x(556) & x(557) & x(582) & x(583) & x(584) & x(610) & x(695) & x(733);
    y(229) <= not(p229_out);
    p229 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110010110000000000000000000011",
            TABLE => "0000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010011000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 3,
            B => -117,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p229_in,
            y(0) => p229_out,
            y(1 to 14 - 1) => dummy229
        );


    p230_in <= x(45) & x(46) & x(50) & x(63) & x(64) & x(66) & x(68) & x(69) & x(70) & x(78) & x(186) & x(210) & x(230) & x(231) & x(232) & x(256) & x(257) & x(284) & x(285) & x(298) & x(299) & x(305) & x(309) & x(310) & x(338) & x(339) & x(349) & x(350) & x(361) & x(366) & x(415) & x(446) & x(474) & x(592) & x(695) & x(720) & x(721) & x(723) & x(732);
    y(230) <= not(p230_out);
    p230 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000000000111111111011110011011000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 3,
            B => -35,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p230_in,
            y(0) => p230_out,
            y(1 to 14 - 1) => dummy230
        );


    p231_in <= x(40) & x(41) & x(46) & x(147) & x(200) & x(276) & x(277) & x(304) & x(305) & x(306) & x(318) & x(319) & x(320) & x(321) & x(361) & x(369) & x(389) & x(390) & x(418) & x(446) & x(454) & x(462) & x(473) & x(474) & x(475) & x(489) & x(490) & x(502) & x(622) & x(623) & x(695) & x(705) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723);
    y(231) <= not(p231_out);
    p231 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00011000000000101111111111111100000000",
            TABLE => "101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 3,
            B => -28,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p231_in,
            y(0) => p231_out,
            y(1 to 14 - 1) => dummy231
        );


    p232_in <= x(44) & x(127) & x(180) & x(181) & x(182) & x(183) & x(205) & x(214) & x(220) & x(234) & x(244) & x(246) & x(247) & x(248) & x(260) & x(275) & x(294) & x(295) & x(306) & x(322) & x(362) & x(370) & x(389) & x(390) & x(396) & x(398) & x(400) & x(418) & x(434) & x(446) & x(462) & x(490) & x(500) & x(528) & x(555) & x(582) & x(657) & x(715) & x(717);
    y(232) <= not(p232_out);
    p232 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111111111100101011000101001111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 2,
            B => 70,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p232_in,
            y(0) => p232_out,
            y(1 to 13 - 1) => dummy232
        );


    p233_in <= x(104) & x(109) & x(122) & x(124) & x(133) & x(134) & x(150) & x(151) & x(212) & x(228) & x(248) & x(249) & x(250) & x(275) & x(276) & x(277) & x(303) & x(304) & x(305) & x(306) & x(333) & x(334) & x(359) & x(360) & x(362) & x(387) & x(388) & x(390) & x(391) & x(418) & x(446) & x(474) & x(502) & x(508) & x(509) & x(526) & x(534) & x(552) & x(554) & x(555) & x(582) & x(584) & x(610) & x(611) & x(638) & x(666) & x(668) & x(696) & x(713) & x(715) & x(716) & x(717) & x(718) & x(720) & x(721) & x(732) & x(733) & x(737) & x(738) & x(739) & x(740) & x(741) & x(742) & x(744) & x(745) & x(746) & x(750);
    y(233) <= not(p233_out);
    p233 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111001110111111111111001001111111110111111111111111111111111111111",
            TABLE => "0000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => 304,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p233_in,
            y(0) => p233_out,
            y(1 to 15 - 1) => dummy233
        );


    p234_in <= x(48) & x(66) & x(117) & x(145) & x(172) & x(219) & x(220) & x(221) & x(228) & x(247) & x(248) & x(249) & x(276) & x(277) & x(305) & x(306) & x(307) & x(325) & x(328) & x(329) & x(330) & x(450) & x(528) & x(583) & x(610) & x(611) & x(687) & x(705) & x(708) & x(720);
    y(234) <= not(p234_out);
    p234 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110001110111111110000011111000",
            TABLE => "010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => 62,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p234_in,
            y(0) => p234_out,
            y(1 to 14 - 1) => dummy234
        );


    p235_in <= x(40) & x(98) & x(181) & x(182) & x(183) & x(184) & x(185) & x(186) & x(213) & x(228) & x(256) & x(276) & x(310) & x(311) & x(338) & x(369) & x(411) & x(438) & x(443) & x(446) & x(462) & x(463) & x(471) & x(473) & x(474) & x(490) & x(491) & x(499) & x(501) & x(518) & x(529) & x(539) & x(540) & x(542) & x(569) & x(719) & x(720) & x(721) & x(732);
    y(235) <= not(p235_out);
    p235 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111001000100100010000100011111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => 2,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p235_in,
            y(0) => p235_out,
            y(1 to 13 - 1) => dummy235
        );


    p236_in <= x(106) & x(198) & x(202) & x(255) & x(256) & x(268) & x(285) & x(294) & x(295) & x(309) & x(310) & x(312) & x(321) & x(322) & x(323) & x(338) & x(339) & x(358) & x(361) & x(362) & x(366) & x(373) & x(391) & x(402) & x(403) & x(418) & x(474) & x(502) & x(557) & x(622) & x(623) & x(677) & x(692) & x(693) & x(694) & x(695) & x(732);
    y(236) <= not(p236_out);
    p236 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000000000000000010001011000000011111",
            TABLE => "1110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101101101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => -95,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p236_in,
            y(0) => p236_out,
            y(1 to 14 - 1) => dummy236
        );


    p237_in <= x(192) & x(193) & x(194) & x(219) & x(220) & x(221) & x(247) & x(248) & x(249) & x(250) & x(256) & x(275) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(320) & x(321) & x(330) & x(333) & x(341) & x(342) & x(347) & x(348) & x(358) & x(359) & x(360) & x(369) & x(370) & x(473) & x(501) & x(515) & x(516) & x(675);
    y(237) <= not(p237_out);
    p237 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000000000100000000001000001110011110",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => -120,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p237_in,
            y(0) => p237_out,
            y(1 to 14 - 1) => dummy237
        );


    p238_in <= x(89) & x(93) & x(94) & x(95) & x(96) & x(97) & x(98) & x(101) & x(118) & x(121) & x(122) & x(123) & x(124) & x(125) & x(126) & x(127) & x(135) & x(149) & x(150) & x(151) & x(152) & x(161) & x(163) & x(189) & x(190) & x(191) & x(355) & x(359) & x(387) & x(390) & x(391) & x(418) & x(473) & x(474) & x(502) & x(520) & x(541) & x(547) & x(548) & x(569) & x(584) & x(720) & x(736) & x(737) & x(738) & x(740) & x(742) & x(745) & x(746) & x(747);
    y(238) <= not(p238_out);
    p238 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111111111110111100000100111111111111111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 2,
            B => 114,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p238_in,
            y(0) => p238_out,
            y(1 to 13 - 1) => dummy238
        );


    p239_in <= x(44) & x(94) & x(95) & x(96) & x(98) & x(118) & x(122) & x(135) & x(163) & x(190) & x(191) & x(192) & x(218) & x(219) & x(220) & x(221) & x(238) & x(247) & x(248) & x(249) & x(254) & x(275) & x(276) & x(277) & x(305) & x(306) & x(328) & x(329) & x(330) & x(331) & x(332) & x(342) & x(358) & x(359) & x(360) & x(361) & x(369) & x(370) & x(388) & x(389) & x(390) & x(391) & x(396) & x(418) & x(446) & x(453) & x(473) & x(474) & x(475) & x(501) & x(502) & x(529) & x(531) & x(619) & x(697) & x(736) & x(738) & x(745) & x(746) & x(747);
    y(239) <= not(p239_out);
    p239 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000011111111101111111110000010000110000100000000000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => -92,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p239_in,
            y(0) => p239_out,
            y(1 to 15 - 1) => dummy239
        );


    p240_in <= x(238) & x(266) & x(267) & x(276) & x(277) & x(304) & x(305) & x(306) & x(344) & x(359) & x(370) & x(387) & x(390) & x(391) & x(397) & x(418) & x(451) & x(473) & x(474) & x(479) & x(502) & x(529) & x(661) & x(720) & x(721) & x(736) & x(737) & x(738) & x(740) & x(741) & x(742) & x(743);
    y(240) <= not(p240_out);
    p240 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111000011011111110111111111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 3,
            B => 151,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p240_in,
            y(0) => p240_out,
            y(1 to 14 - 1) => dummy240
        );


    p241_in <= x(35) & x(108) & x(192) & x(248) & x(249) & x(276) & x(277) & x(305) & x(330) & x(331) & x(332) & x(334) & x(358) & x(359) & x(360) & x(379) & x(387) & x(388) & x(389) & x(407) & x(416) & x(418) & x(425) & x(454) & x(473) & x(501) & x(519) & x(520) & x(528) & x(529) & x(544) & x(545) & x(546) & x(569) & x(571) & x(572) & x(573) & x(697);
    y(241) <= not(p241_out);
    p241 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11000000111011101110111111111111111111",
            TABLE => "100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 2,
            B => 58,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p241_in,
            y(0) => p241_out,
            y(1 to 13 - 1) => dummy241
        );


    p242_in <= x(209) & x(210) & x(211) & x(238) & x(247) & x(248) & x(256) & x(275) & x(276) & x(277) & x(303) & x(304) & x(305) & x(306) & x(332) & x(333) & x(415) & x(443) & x(444) & x(462) & x(489) & x(490) & x(636) & x(663) & x(697) & x(705) & x(718) & x(719) & x(721) & x(722) & x(747);
    y(242) <= not(p242_out);
    p242 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111110111111111111000000111111",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 3,
            B => 75,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p242_in,
            y(0) => p242_out,
            y(1 to 14 - 1) => dummy242
        );


    p243_in <= x(192) & x(220) & x(221) & x(248) & x(249) & x(276) & x(277) & x(304) & x(305) & x(306) & x(320) & x(329) & x(330) & x(331) & x(346) & x(347) & x(348) & x(356) & x(357) & x(358) & x(360) & x(369) & x(389) & x(391) & x(418) & x(443) & x(473) & x(474) & x(502) & x(514) & x(515) & x(516) & x(517) & x(675) & x(676) & x(679) & x(697) & x(705) & x(706) & x(708) & x(711) & x(722);
    y(243) <= not(p243_out);
    p243 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111111110001110000100010000000111011111",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => 42,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p243_in,
            y(0) => p243_out,
            y(1 to 14 - 1) => dummy243
        );


    p244_in <= x(44) & x(89) & x(135) & x(162) & x(163) & x(184) & x(191) & x(211) & x(212) & x(213) & x(238) & x(239) & x(240) & x(250) & x(303) & x(304) & x(310) & x(331) & x(332) & x(338) & x(339) & x(366) & x(411) & x(438) & x(471) & x(489) & x(490) & x(499) & x(517) & x(518) & x(611) & x(720) & x(747);
    y(244) <= not(p244_out);
    p244 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001110100000000010011111011011100",
            TABLE => "001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001100011101001011011111111",
            SHIFT => 2,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p244_in,
            y(0) => p244_out,
            y(1 to 13 - 1) => dummy244
        );


    p245_in <= x(44) & x(96) & x(97) & x(98) & x(99) & x(171) & x(199) & x(219) & x(220) & x(248) & x(255) & x(266) & x(267) & x(275) & x(276) & x(283) & x(294) & x(295) & x(296) & x(309) & x(310) & x(321) & x(322) & x(323) & x(338) & x(339) & x(340) & x(362) & x(366) & x(375) & x(391) & x(398) & x(399) & x(403) & x(418) & x(427) & x(428) & x(431) & x(637) & x(663) & x(664) & x(665) & x(677) & x(705) & x(707) & x(708) & x(709) & x(710) & x(711) & x(712) & x(713) & x(714) & x(715) & x(716) & x(717) & x(718) & x(719) & x(720) & x(721) & x(736) & x(737) & x(738) & x(739) & x(741) & x(742) & x(743) & x(744) & x(745) & x(746) & x(747) & x(748) & x(750) & x(764) & x(774);
    y(245) <= not(p245_out);
    p245 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000001110001100000000000000101110111111100000000000000000000000000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 2,
            B => -156,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p245_in,
            y(0) => p245_out,
            y(1 to 14 - 1) => dummy245
        );


    p246_in <= x(104) & x(105) & x(106) & x(134) & x(135) & x(162) & x(163) & x(222) & x(305) & x(321) & x(330) & x(331) & x(332) & x(359) & x(360) & x(717) & x(720);
    y(246) <= not(p246_out);
    p246 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111100000000",
            TABLE => "00000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100100000000100000001000000011101000100000001110100011101000111111100001011110000001100000011110100010000001111010001110100001111110011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 54,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p246_in,
            y(0) => p246_out,
            y(1 to 14 - 1) => dummy246
        );


    p247_in <= x(73) & x(145) & x(161) & x(247) & x(248) & x(276) & x(277) & x(309) & x(338) & x(348) & x(366) & x(375) & x(380) & x(388) & x(398) & x(400) & x(401) & x(437) & x(450) & x(464) & x(465) & x(492) & x(493) & x(507) & x(520) & x(535) & x(542) & x(544) & x(694) & x(705) & x(739) & x(743) & x(745);
    y(247) <= not(p247_out);
    p247 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010000000101111111111111110011000",
            TABLE => "111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 2,
            B => -29,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p247_in,
            y(0) => p247_out,
            y(1 to 13 - 1) => dummy247
        );


    p248_in <= x(70) & x(91) & x(106) & x(108) & x(146) & x(165) & x(187) & x(188) & x(189) & x(190) & x(191) & x(192) & x(216) & x(217) & x(218) & x(219) & x(220) & x(242) & x(243) & x(244) & x(245) & x(246) & x(247) & x(248) & x(249) & x(272) & x(273) & x(274) & x(275) & x(276) & x(277) & x(278) & x(292) & x(305) & x(306) & x(307) & x(334) & x(378) & x(390) & x(426) & x(490) & x(500) & x(537) & x(545) & x(573) & x(574) & x(656) & x(657) & x(658) & x(659) & x(683) & x(687) & x(688) & x(705) & x(733) & x(734) & x(735) & x(736) & x(737) & x(738) & x(740) & x(741) & x(742) & x(746);
    y(248) <= not(p248_out);
    p248 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111100000000000000000000000000000000101100111000000011111111111",
            TABLE => "0000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101100000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101101111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 2,
            B => -32,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p248_in,
            y(0) => p248_out,
            y(1 to 14 - 1) => dummy248
        );


    p249_in <= x(46) & x(65) & x(101) & x(156) & x(204) & x(205) & x(220) & x(221) & x(231) & x(248) & x(249) & x(259) & x(260) & x(275) & x(276) & x(277) & x(286) & x(305) & x(306) & x(307) & x(313) & x(314) & x(330) & x(334) & x(350) & x(358) & x(359) & x(361) & x(389) & x(390) & x(391) & x(418) & x(446) & x(473) & x(500) & x(501) & x(527) & x(528) & x(556) & x(582) & x(583) & x(609) & x(610) & x(611) & x(631) & x(634) & x(635) & x(636) & x(637) & x(638) & x(658) & x(659) & x(660) & x(661) & x(662) & x(663) & x(664) & x(665) & x(688) & x(695) & x(705) & x(720) & x(721) & x(723) & x(732) & x(733) & x(769);
    y(249) <= not(p249_out);
    p249 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0101111111111111111111010001111111111111111111111111111111100000001",
            TABLE => "0001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 2,
            B => 132,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p249_in,
            y(0) => p249_out,
            y(1 to 14 - 1) => dummy249
        );


    p250_in <= x(118) & x(144) & x(145) & x(171) & x(172) & x(174) & x(192) & x(199) & x(200) & x(201) & x(220) & x(227) & x(228) & x(248) & x(249) & x(255) & x(256) & x(275) & x(276) & x(277) & x(283) & x(290) & x(296) & x(299) & x(305) & x(306) & x(310) & x(311) & x(329) & x(330) & x(331) & x(334) & x(338) & x(339) & x(359) & x(360) & x(366) & x(375) & x(376) & x(388) & x(403) & x(405) & x(407) & x(411) & x(422) & x(438) & x(439) & x(466) & x(467) & x(474) & x(493) & x(500) & x(502) & x(530) & x(535) & x(557) & x(558) & x(563) & x(564) & x(648) & x(649) & x(650) & x(676) & x(677) & x(678) & x(690) & x(692) & x(695) & x(704) & x(705) & x(706) & x(707) & x(708) & x(709) & x(774);
    y(250) <= not(p250_out);
    p250 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000100010011001110100110000010000011011100000000100000000000001110000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 2,
            B => -176,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p250_in,
            y(0) => p250_out,
            y(1 to 14 - 1) => dummy250
        );


    p251_in <= x(210) & x(271) & x(305) & x(322) & x(323) & x(330) & x(331) & x(332) & x(350) & x(351) & x(358) & x(359) & x(360) & x(361) & x(368) & x(378) & x(387) & x(388) & x(389) & x(390) & x(405) & x(406) & x(407) & x(474) & x(500) & x(527) & x(528) & x(578) & x(603) & x(604) & x(605) & x(606) & x(695) & x(705) & x(707) & x(709) & x(718) & x(719) & x(720) & x(721) & x(722) & x(723) & x(745) & x(746);
    y(251) <= not(p251_out);
    p251 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01000111001111001111000111111111000000000000",
            TABLE => "110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 2,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p251_in,
            y(0) => p251_out,
            y(1 to 13 - 1) => dummy251
        );


    p252_in <= x(192) & x(220) & x(221) & x(248) & x(249) & x(276) & x(277) & x(304) & x(305) & x(306) & x(329) & x(330) & x(331) & x(333) & x(358) & x(359) & x(360) & x(366) & x(386) & x(387) & x(388) & x(391) & x(416) & x(418) & x(424) & x(455) & x(474) & x(485) & x(529) & x(717) & x(718) & x(737) & x(739) & x(743) & x(744) & x(745) & x(746) & x(747) & x(750);
    y(252) <= not(p252_out);
    p252 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000000011101110111010110100000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 3,
            B => -104,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p252_in,
            y(0) => p252_out,
            y(1 to 14 - 1) => dummy252
        );


    p253_in <= x(41) & x(96) & x(97) & x(98) & x(99) & x(100) & x(101) & x(145) & x(161) & x(162) & x(163) & x(165) & x(171) & x(190) & x(191) & x(192) & x(199) & x(218) & x(219) & x(220) & x(221) & x(248) & x(249) & x(260) & x(276) & x(277) & x(289) & x(290) & x(291) & x(305) & x(306) & x(307) & x(325) & x(326) & x(327) & x(328) & x(329) & x(330) & x(334) & x(354) & x(376) & x(390) & x(528) & x(583) & x(610) & x(611) & x(637) & x(657) & x(663) & x(664) & x(665) & x(676) & x(697) & x(705) & x(707) & x(708) & x(709) & x(719) & x(720) & x(721) & x(735) & x(736) & x(742) & x(745) & x(746) & x(747);
    y(253) <= not(p253_out);
    p253 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000001111011101111111111111110000001011111111111010000000000000",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 2,
            B => 17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p253_in,
            y(0) => p253_out,
            y(1 to 14 - 1) => dummy253
        );


    p254_in <= x(70) & x(71) & x(72) & x(108) & x(145) & x(248) & x(249) & x(250) & x(277) & x(305) & x(306) & x(321) & x(322) & x(323) & x(333) & x(343) & x(387) & x(426) & x(453) & x(454) & x(481) & x(482) & x(501) & x(509) & x(510) & x(511) & x(528) & x(538) & x(545) & x(565) & x(657) & x(718) & x(719) & x(774);
    y(254) <= not(p254_out);
    p254 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110111111111111000000000000001111",
            TABLE => "0000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 2,
            B => 16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p254_in,
            y(0) => p254_out,
            y(1 to 13 - 1) => dummy254
        );


    p255_in <= x(106) & x(192) & x(193) & x(217) & x(218) & x(219) & x(220) & x(221) & x(242) & x(243) & x(244) & x(247) & x(248) & x(249) & x(250) & x(274) & x(275) & x(276) & x(277) & x(278) & x(303) & x(304) & x(305) & x(306) & x(333) & x(334) & x(390) & x(470) & x(510) & x(540) & x(552) & x(568) & x(571) & x(580) & x(592) & x(597) & x(625) & x(647);
    y(255) <= not(p255_out);
    p255 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000000000000000000000000000000000000",
            TABLE => "111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 2,
            B => -135,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p255_in,
            y(0) => p255_out,
            y(1 to 13 - 1) => dummy255
        );



--    p1 : perceptron
--        Generic map (
--            WEIGHTS => "",
--            SHIFT => "",
--            B => "",
--            BATCH_POSITIVE => ""
--        )
--        Port map (
--            x => x(0) & x(2) & ...,
--            y => ""
--        );

end layer_1;

architecture layer_2 of layer is

    Component perceptron
    Generic (
        WEIGHTS : STD_LOGIC_VECTOR;
        SHIFT : Integer;     -- number of shift (left + or right -)
        B : Integer;          -- bias of batch norm
        BATCH_POSITIVE : Boolean    
    );
    Port ( 
        x : in STD_LOGIC_VECTOR;
        y : out STD_LOGIC_VECTOR
   );
    end component;
    
    -- Signals
    signal p0_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p0_out : STD_LOGIC;
	signal p1_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p1_out : STD_LOGIC;
	signal p2_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p2_out : STD_LOGIC;
	signal p3_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p3_out : STD_LOGIC;
	signal p4_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p4_out : STD_LOGIC;
	signal p5_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p5_out : STD_LOGIC;
	signal p6_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p6_out : STD_LOGIC;
	signal p7_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p7_out : STD_LOGIC;
	signal p8_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p8_out : STD_LOGIC;
	signal p9_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p9_out : STD_LOGIC;
	signal p10_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p10_out : STD_LOGIC;
	signal p11_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p11_out : STD_LOGIC;
	signal p12_in : STD_LOGIC_VECTOR(0 to 45 - 1);
	signal p12_out : STD_LOGIC;
	signal p13_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p13_out : STD_LOGIC;
	signal p14_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p14_out : STD_LOGIC;
	signal p15_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p15_out : STD_LOGIC;
	signal p16_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p16_out : STD_LOGIC;
	signal p17_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p17_out : STD_LOGIC;
	signal p18_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p18_out : STD_LOGIC;
	signal p19_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p19_out : STD_LOGIC;
	signal p20_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p20_out : STD_LOGIC;
	signal p21_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p21_out : STD_LOGIC;
	signal p22_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p22_out : STD_LOGIC;
	signal p23_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p23_out : STD_LOGIC;
	signal p24_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p24_out : STD_LOGIC;
	signal p25_in : STD_LOGIC_VECTOR(0 to 52 - 1);
	signal p25_out : STD_LOGIC;
	signal p26_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p26_out : STD_LOGIC;
	signal p27_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p27_out : STD_LOGIC;
	signal p28_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p28_out : STD_LOGIC;
	signal p29_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p29_out : STD_LOGIC;
	signal p30_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p30_out : STD_LOGIC;
	signal p31_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p31_out : STD_LOGIC;
	signal p32_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p32_out : STD_LOGIC;
	signal p33_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p33_out : STD_LOGIC;
	signal p34_in : STD_LOGIC_VECTOR(0 to 46 - 1);
	signal p34_out : STD_LOGIC;
	signal p35_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p35_out : STD_LOGIC;
	signal p36_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p36_out : STD_LOGIC;
	signal p37_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p37_out : STD_LOGIC;
	signal p38_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p38_out : STD_LOGIC;
	signal p39_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p39_out : STD_LOGIC;
	signal p40_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p40_out : STD_LOGIC;
	signal p41_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p41_out : STD_LOGIC;
	signal p42_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p42_out : STD_LOGIC;
	signal p43_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p43_out : STD_LOGIC;
	signal p44_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p44_out : STD_LOGIC;
	signal p45_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p45_out : STD_LOGIC;
	signal p46_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p46_out : STD_LOGIC;
	signal p47_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p47_out : STD_LOGIC;
	signal p48_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p48_out : STD_LOGIC;
	signal p49_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p49_out : STD_LOGIC;
	signal p50_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p50_out : STD_LOGIC;
	signal p51_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p51_out : STD_LOGIC;
	signal p52_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p52_out : STD_LOGIC;
	signal p53_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p53_out : STD_LOGIC;
	signal p54_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p54_out : STD_LOGIC;
	signal p55_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p55_out : STD_LOGIC;
	signal p56_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p56_out : STD_LOGIC;
	signal p57_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p57_out : STD_LOGIC;
	signal p58_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p58_out : STD_LOGIC;
	signal p59_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p59_out : STD_LOGIC;
	signal p60_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p60_out : STD_LOGIC;
	signal p61_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p61_out : STD_LOGIC;
	signal p62_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p62_out : STD_LOGIC;
	signal p63_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p63_out : STD_LOGIC;
	signal p64_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p64_out : STD_LOGIC;
	signal p65_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p65_out : STD_LOGIC;
	signal p66_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p66_out : STD_LOGIC;
	signal p67_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p67_out : STD_LOGIC;
	signal p68_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p68_out : STD_LOGIC;
	signal p69_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p69_out : STD_LOGIC;
	signal p70_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p70_out : STD_LOGIC;
	signal p71_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p71_out : STD_LOGIC;
	signal p72_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p72_out : STD_LOGIC;
	signal p73_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p73_out : STD_LOGIC;
	signal p74_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p74_out : STD_LOGIC;
	signal p75_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p75_out : STD_LOGIC;
	signal p76_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p76_out : STD_LOGIC;
	signal p77_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p77_out : STD_LOGIC;
	signal p78_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p78_out : STD_LOGIC;
	signal p79_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p79_out : STD_LOGIC;
	signal p80_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p80_out : STD_LOGIC;
	signal p81_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p81_out : STD_LOGIC;
	signal p82_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p82_out : STD_LOGIC;
	signal p83_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p83_out : STD_LOGIC;
	signal p84_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p84_out : STD_LOGIC;
	signal p85_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p85_out : STD_LOGIC;
	signal p86_in : STD_LOGIC_VECTOR(0 to 48 - 1);
	signal p86_out : STD_LOGIC;
	signal p87_in : STD_LOGIC_VECTOR(0 to 48 - 1);
	signal p87_out : STD_LOGIC;
	signal p88_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p88_out : STD_LOGIC;
	signal p89_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p89_out : STD_LOGIC;
	signal p90_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p90_out : STD_LOGIC;
	signal p91_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p91_out : STD_LOGIC;
	signal p92_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p92_out : STD_LOGIC;
	signal p93_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p93_out : STD_LOGIC;
	signal p94_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p94_out : STD_LOGIC;
	signal p95_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p95_out : STD_LOGIC;
	signal p96_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p96_out : STD_LOGIC;
	signal p97_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p97_out : STD_LOGIC;
	signal p98_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p98_out : STD_LOGIC;
	signal p99_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p99_out : STD_LOGIC;
	signal p100_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p100_out : STD_LOGIC;
	signal p101_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p101_out : STD_LOGIC;
	signal p102_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p102_out : STD_LOGIC;
	signal p103_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p103_out : STD_LOGIC;
	signal p104_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p104_out : STD_LOGIC;
	signal p105_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p105_out : STD_LOGIC;
	signal p106_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p106_out : STD_LOGIC;
	signal p107_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p107_out : STD_LOGIC;
	signal p108_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p108_out : STD_LOGIC;
	signal p109_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p109_out : STD_LOGIC;
	signal p110_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p110_out : STD_LOGIC;
	signal p111_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p111_out : STD_LOGIC;
	signal p112_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p112_out : STD_LOGIC;
	signal p113_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p113_out : STD_LOGIC;
	signal p114_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p114_out : STD_LOGIC;
	signal p115_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p115_out : STD_LOGIC;
	signal p116_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p116_out : STD_LOGIC;
	signal p117_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p117_out : STD_LOGIC;
	signal p118_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p118_out : STD_LOGIC;
	signal p119_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p119_out : STD_LOGIC;
	signal p120_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p120_out : STD_LOGIC;
	signal p121_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p121_out : STD_LOGIC;
	signal p122_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p122_out : STD_LOGIC;
	signal p123_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p123_out : STD_LOGIC;
	signal p124_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p124_out : STD_LOGIC;
	signal p125_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p125_out : STD_LOGIC;
	signal p126_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p126_out : STD_LOGIC;
	signal p127_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p127_out : STD_LOGIC;
	signal p128_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p128_out : STD_LOGIC;
	signal p129_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p129_out : STD_LOGIC;
	signal p130_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p130_out : STD_LOGIC;
	signal p131_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p131_out : STD_LOGIC;
	signal p132_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p132_out : STD_LOGIC;
	signal p133_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p133_out : STD_LOGIC;
	signal p134_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p134_out : STD_LOGIC;
	signal p135_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p135_out : STD_LOGIC;
	signal p136_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p136_out : STD_LOGIC;
	signal p137_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p137_out : STD_LOGIC;
	signal p138_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p138_out : STD_LOGIC;
	signal p139_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p139_out : STD_LOGIC;
	signal p140_in : STD_LOGIC_VECTOR(0 to 45 - 1);
	signal p140_out : STD_LOGIC;
	signal p141_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p141_out : STD_LOGIC;
	signal p142_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p142_out : STD_LOGIC;
	signal p143_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p143_out : STD_LOGIC;
	signal p144_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p144_out : STD_LOGIC;
	signal p145_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p145_out : STD_LOGIC;
	signal p146_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p146_out : STD_LOGIC;
	signal p147_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p147_out : STD_LOGIC;
	signal p148_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p148_out : STD_LOGIC;
	signal p149_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p149_out : STD_LOGIC;
	signal p150_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p150_out : STD_LOGIC;
	signal p151_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p151_out : STD_LOGIC;
	signal p152_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p152_out : STD_LOGIC;
	signal p153_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p153_out : STD_LOGIC;
	signal p154_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p154_out : STD_LOGIC;
	signal p155_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p155_out : STD_LOGIC;
	signal p156_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p156_out : STD_LOGIC;
	signal p157_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p157_out : STD_LOGIC;
	signal p158_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p158_out : STD_LOGIC;
	signal p159_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p159_out : STD_LOGIC;
	signal p160_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p160_out : STD_LOGIC;
	signal p161_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p161_out : STD_LOGIC;
	signal p162_in : STD_LOGIC_VECTOR(0 to 44 - 1);
	signal p162_out : STD_LOGIC;
	signal p163_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p163_out : STD_LOGIC;
	signal p164_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p164_out : STD_LOGIC;
	signal p165_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p165_out : STD_LOGIC;
	signal p166_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p166_out : STD_LOGIC;
	signal p167_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p167_out : STD_LOGIC;
	signal p168_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p168_out : STD_LOGIC;
	signal p169_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p169_out : STD_LOGIC;
	signal p170_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p170_out : STD_LOGIC;
	signal p171_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p171_out : STD_LOGIC;
	signal p172_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p172_out : STD_LOGIC;
	signal p173_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p173_out : STD_LOGIC;
	signal p174_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p174_out : STD_LOGIC;
	signal p175_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p175_out : STD_LOGIC;
	signal p176_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p176_out : STD_LOGIC;
	signal p177_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p177_out : STD_LOGIC;
	signal p178_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p178_out : STD_LOGIC;
	signal p179_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p179_out : STD_LOGIC;
	signal p180_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p180_out : STD_LOGIC;
	signal p181_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p181_out : STD_LOGIC;
	signal p182_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p182_out : STD_LOGIC;
	signal p183_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p183_out : STD_LOGIC;
	signal p184_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p184_out : STD_LOGIC;
	signal p185_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p185_out : STD_LOGIC;
	signal p186_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p186_out : STD_LOGIC;
	signal p187_in : STD_LOGIC_VECTOR(0 to 49 - 1);
	signal p187_out : STD_LOGIC;
	signal p188_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p188_out : STD_LOGIC;
	signal p189_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p189_out : STD_LOGIC;
	signal p190_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p190_out : STD_LOGIC;
	signal p191_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p191_out : STD_LOGIC;
	signal p192_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p192_out : STD_LOGIC;
	signal p193_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p193_out : STD_LOGIC;
	signal p194_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p194_out : STD_LOGIC;
	signal p195_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p195_out : STD_LOGIC;
	signal p196_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p196_out : STD_LOGIC;
	signal p197_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p197_out : STD_LOGIC;
	signal p198_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p198_out : STD_LOGIC;
	signal p199_in : STD_LOGIC_VECTOR(0 to 47 - 1);
	signal p199_out : STD_LOGIC;
	signal p200_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p200_out : STD_LOGIC;
	signal p201_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p201_out : STD_LOGIC;
	signal p202_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p202_out : STD_LOGIC;
	signal p203_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p203_out : STD_LOGIC;
	signal p204_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p204_out : STD_LOGIC;
	signal p205_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p205_out : STD_LOGIC;
	signal p206_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p206_out : STD_LOGIC;
	signal p207_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p207_out : STD_LOGIC;
	signal p208_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p208_out : STD_LOGIC;
	signal p209_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p209_out : STD_LOGIC;
	signal p210_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p210_out : STD_LOGIC;
	signal p211_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p211_out : STD_LOGIC;
	signal p212_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p212_out : STD_LOGIC;
	signal p213_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p213_out : STD_LOGIC;
	signal p214_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p214_out : STD_LOGIC;
	signal p215_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p215_out : STD_LOGIC;
	signal p216_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p216_out : STD_LOGIC;
	signal p217_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p217_out : STD_LOGIC;
	signal p218_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p218_out : STD_LOGIC;
	signal p219_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p219_out : STD_LOGIC;
	signal p220_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p220_out : STD_LOGIC;
	signal p221_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p221_out : STD_LOGIC;
	signal p222_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p222_out : STD_LOGIC;
	signal p223_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p223_out : STD_LOGIC;
	signal p224_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p224_out : STD_LOGIC;
	signal p225_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p225_out : STD_LOGIC;
	signal p226_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p226_out : STD_LOGIC;
	signal p227_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p227_out : STD_LOGIC;
	signal p228_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p228_out : STD_LOGIC;
	signal p229_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p229_out : STD_LOGIC;
	signal p230_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p230_out : STD_LOGIC;
	signal p231_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p231_out : STD_LOGIC;
	signal p232_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p232_out : STD_LOGIC;
	signal p233_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p233_out : STD_LOGIC;
	signal p234_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p234_out : STD_LOGIC;
	signal p235_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p235_out : STD_LOGIC;
	signal p236_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p236_out : STD_LOGIC;
	signal p237_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p237_out : STD_LOGIC;
	signal p238_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p238_out : STD_LOGIC;
	signal p239_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p239_out : STD_LOGIC;
	signal p240_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p240_out : STD_LOGIC;
	signal p241_in : STD_LOGIC_VECTOR(0 to 44 - 1);
	signal p241_out : STD_LOGIC;
	signal p242_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p242_out : STD_LOGIC;
	signal p243_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p243_out : STD_LOGIC;
	signal p244_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p244_out : STD_LOGIC;
	signal p245_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p245_out : STD_LOGIC;
	signal p246_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p246_out : STD_LOGIC;
	signal p247_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p247_out : STD_LOGIC;
	signal p248_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p248_out : STD_LOGIC;
	signal p249_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p249_out : STD_LOGIC;
	signal p250_in : STD_LOGIC_VECTOR(0 to 49 - 1);
	signal p250_out : STD_LOGIC;
	signal p251_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p251_out : STD_LOGIC;
	signal p252_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p252_out : STD_LOGIC;
	signal p253_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p253_out : STD_LOGIC;
	signal p254_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p254_out : STD_LOGIC;
	signal p255_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p255_out : STD_LOGIC;
	
    
    -- Dummies
    signal dummy0 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy1 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy2 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy3 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy4 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy5 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy6 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy7 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy8 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy9 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy10 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy11 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy12 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy13 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy14 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy15 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy16 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy17 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy18 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy19 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy20 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy21 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy22 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy23 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy24 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy25 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy26 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy27 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy28 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy29 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy30 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy31 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy32 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy33 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy34 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy35 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy36 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy37 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy38 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy39 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy40 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy41 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy42 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy43 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy44 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy45 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy46 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy47 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy48 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy49 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy50 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy51 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy52 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy53 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy54 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy55 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy56 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy57 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy58 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy59 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy60 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy61 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy62 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy63 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy64 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy65 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy66 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy67 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy68 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy69 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy70 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy71 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy72 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy73 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy74 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy75 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy76 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy77 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy78 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy79 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy80 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy81 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy82 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy83 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy84 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy85 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy86 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy87 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy88 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy89 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy90 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy91 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy92 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy93 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy94 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy95 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy96 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy97 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy98 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy99 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy100 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy101 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy102 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy103 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy104 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy105 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy106 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy107 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy108 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy109 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy110 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy111 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy112 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy113 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy114 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy115 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy116 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy117 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy118 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy119 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy120 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy121 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy122 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy123 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy124 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy125 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy126 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy127 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy128 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy129 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy130 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy131 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy132 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy133 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy134 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy135 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy136 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy137 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy138 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy139 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy140 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy141 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy142 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy143 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy144 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy145 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy146 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy147 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy148 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy149 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy150 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy151 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy152 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy153 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy154 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy155 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy156 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy157 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy158 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy159 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy160 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy161 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy162 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy163 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy164 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy165 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy166 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy167 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy168 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy169 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy170 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy171 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy172 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy173 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy174 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy175 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy176 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy177 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy178 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy179 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy180 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy181 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy182 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy183 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy184 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy185 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy186 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy187 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy188 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy189 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy190 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy191 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy192 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy193 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy194 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy195 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy196 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy197 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy198 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy199 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy200 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy201 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy202 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy203 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy204 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy205 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy206 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy207 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy208 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy209 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy210 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy211 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy212 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy213 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy214 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy215 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy216 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy217 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy218 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy219 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy220 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy221 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy222 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy223 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy224 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy225 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy226 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy227 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy228 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy229 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy230 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy231 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy232 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy233 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy234 : STD_LOGIC_VECTOR(0 to 16 - 2);
	signal dummy235 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy236 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy237 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy238 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy239 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy240 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy241 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy242 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy243 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy244 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy245 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy246 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy247 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy248 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy249 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy250 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy251 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy252 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy253 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy254 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy255 : STD_LOGIC_VECTOR(0 to 15 - 2);
	 
    
begin

    
    p0_in <= x(11) & x(16) & x(19) & x(27) & x(28) & x(38) & x(48) & x(49) & x(50) & x(53) & x(56) & x(61) & x(65) & x(77) & x(89) & x(107) & x(126) & x(139) & x(145) & x(150) & x(151) & x(156) & x(175) & x(177) & x(189) & x(210) & x(218) & x(232);
    y(0) <= not(p0_out);
    p0 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000001100011101000110111010",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101100000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101100001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010010000010110010001001001011001001101001100101100000000000000000",
            SHIFT => 4,
            B => -19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p0_in,
            y(0) => p0_out,
            y(1 to 14 - 1) => dummy0
        );


    p1_in <= x(6) & x(10) & x(24) & x(33) & x(47) & x(54) & x(61) & x(66) & x(70) & x(72) & x(74) & x(79) & x(88) & x(89) & x(96) & x(97) & x(99) & x(101) & x(108) & x(121) & x(122) & x(127) & x(135) & x(144) & x(161) & x(175) & x(177) & x(184) & x(211) & x(212) & x(216) & x(220) & x(231) & x(232) & x(234) & x(242) & x(248) & x(249) & x(253);
    y(1) <= not(p1_out);
    p1 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111000000001001101100110110100111010111",
            TABLE => "000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 4,
            B => 43,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p1_in,
            y(0) => p1_out,
            y(1 to 15 - 1) => dummy1
        );


    p2_in <= x(4) & x(5) & x(10) & x(13) & x(18) & x(22) & x(25) & x(32) & x(52) & x(69) & x(72) & x(74) & x(79) & x(87) & x(91) & x(92) & x(93) & x(94) & x(98) & x(142) & x(143) & x(154) & x(167) & x(171) & x(172) & x(179) & x(181) & x(189) & x(196) & x(206) & x(210) & x(225) & x(238) & x(248) & x(249);
    y(2) <= not(p2_out);
    p2 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00100111110010110101110011001100011",
            TABLE => "11010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100100000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100100000100010011010000000000000100010011011101111100000100010011010010010001001101101100100010010001001101110110110010010001001101100101100110100101101001100101100110100110010110100101100110100100001000100011101000111011101111000000000000100000001000100011100001100010001110100011101110011101110001000110000001100010001110011010011001011010010110011010011001011001101001011010011001011000010000000000000111000100010000011100010001000011110111011100010001100010001110011100010001100001110001000110001110011101110001100101100110100101101001100101100110100110010110100101100110100111110111011100010111000100010000111001110111000101110001000110001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p2_in,
            y(0) => p2_out,
            y(1 to 15 - 1) => dummy2
        );


    p3_in <= x(25) & x(27) & x(43) & x(50) & x(74) & x(83) & x(88) & x(98) & x(120) & x(132) & x(134) & x(136) & x(142) & x(153) & x(157) & x(158) & x(167) & x(170) & x(176) & x(177) & x(193) & x(198) & x(199) & x(210) & x(214) & x(218) & x(221) & x(222) & x(236) & x(240) & x(252) & x(254);
    y(3) <= not(p3_out);
    p3 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10001100111111000011010011010101",
            TABLE => "011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 4,
            B => -48,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p3_in,
            y(0) => p3_out,
            y(1 to 15 - 1) => dummy3
        );


    p4_in <= x(0) & x(6) & x(10) & x(20) & x(22) & x(25) & x(27) & x(28) & x(38) & x(39) & x(49) & x(52) & x(65) & x(77) & x(80) & x(87) & x(91) & x(95) & x(113) & x(114) & x(129) & x(142) & x(149) & x(154) & x(156) & x(162) & x(167) & x(169) & x(176) & x(179) & x(185) & x(189) & x(194) & x(197) & x(198) & x(211) & x(230) & x(235) & x(238) & x(242) & x(244);
    y(4) <= not(p4_out);
    p4 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01000000010011010101101001100011110001110",
            TABLE => "11101000100000001111111011101000100000000000000011101000100000001110100010000001011111101110100010000001000101111110100010000001011010011001011010010110011010011001011001101001011010011001011011101111100011101000111000001000100011100000100000001000000000001110011110001110100011100001100010001110000110000001100001110001011010011001011010010110011010011001011001101001011010011001011000000100000000000100110100000100010011010000010011011111010011010010010010110010010011010010010001001101001001001101101101001101100101100110100101101001100101100110100110010110100101100110100100100000101100101011001011111011000000000010000000100000101100100010010010110010101100101101101101001101001001000010010010110010011010011001011010010110011010011001011001101001011010011001011010000000111010001110100011111110000000001000000010000000111010001000000111101000111010000111111000010111100000011000000111101000100101100110100101101001100101100110100110010110100101100110100100000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100100101011101111110000001000101011001010111011110101000010001010110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 28,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p4_in,
            y(0) => p4_out,
            y(1 to 15 - 1) => dummy4
        );


    p5_in <= x(1) & x(7) & x(12) & x(17) & x(56) & x(59) & x(93) & x(119) & x(120) & x(121) & x(127) & x(133) & x(155) & x(156) & x(167) & x(174) & x(175) & x(176) & x(180) & x(189) & x(200) & x(210) & x(212) & x(225) & x(231) & x(232);
    y(5) <= not(p5_out);
    p5 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11110000110010001011100010",
            TABLE => "000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 4,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p5_in,
            y(0) => p5_out,
            y(1 to 14 - 1) => dummy5
        );


    p6_in <= x(0) & x(2) & x(5) & x(10) & x(17) & x(21) & x(23) & x(25) & x(27) & x(35) & x(71) & x(77) & x(80) & x(82) & x(84) & x(88) & x(91) & x(95) & x(96) & x(101) & x(102) & x(110) & x(154) & x(155) & x(156) & x(161) & x(167) & x(179) & x(196) & x(197) & x(208) & x(227) & x(230) & x(233) & x(235) & x(238) & x(242);
    y(6) <= not(p6_out);
    p6 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000000110001001100110111001100010000",
            TABLE => "1110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101101110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p6_in,
            y(0) => p6_out,
            y(1 to 15 - 1) => dummy6
        );


    p7_in <= x(1) & x(7) & x(10) & x(12) & x(25) & x(27) & x(33) & x(34) & x(37) & x(44) & x(50) & x(51) & x(53) & x(62) & x(68) & x(71) & x(87) & x(88) & x(98) & x(119) & x(120) & x(124) & x(127) & x(137) & x(143) & x(148) & x(162) & x(167) & x(172) & x(173) & x(174) & x(198) & x(201) & x(203) & x(209) & x(218) & x(219) & x(227) & x(228) & x(231) & x(232) & x(247) & x(253);
    y(7) <= not(p7_out);
    p7 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111110110010101001011011100110100111101011",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101101000111000001000111011111000111000001000000000001000111000001000100011100001100011100111100011100001100001110001100011100001100010010110011010010110100110010110011010011001011010010110011010010000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010010111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101100000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p7_in,
            y(0) => p7_out,
            y(1 to 15 - 1) => dummy7
        );


    p8_in <= x(2) & x(7) & x(10) & x(33) & x(48) & x(49) & x(53) & x(54) & x(65) & x(71) & x(72) & x(91) & x(96) & x(101) & x(105) & x(106) & x(114) & x(119) & x(133) & x(148) & x(150) & x(156) & x(158) & x(162) & x(167) & x(170) & x(174) & x(175) & x(179) & x(203) & x(206) & x(213) & x(225) & x(230) & x(235) & x(244) & x(249);
    y(8) <= not(p8_out);
    p8 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110010100010101001111000101101111011",
            TABLE => "0100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101101101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010011000111000001000111011111000111000001000000000001000111000001000100011100001100011100111100011100001100001110001100011100001100010010110011010010110100110010110011010011001011010010110011010010000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101100000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p8_in,
            y(0) => p8_out,
            y(1 to 15 - 1) => dummy8
        );


    p9_in <= x(1) & x(13) & x(27) & x(31) & x(35) & x(40) & x(61) & x(69) & x(70) & x(75) & x(80) & x(83) & x(84) & x(85) & x(93) & x(103) & x(104) & x(109) & x(111) & x(113) & x(131) & x(132) & x(139) & x(142) & x(156) & x(161) & x(166) & x(168) & x(177) & x(184) & x(191) & x(193) & x(194) & x(203) & x(205) & x(211) & x(228) & x(233) & x(237) & x(238) & x(242) & x(244) & x(248);
    y(9) <= not(p9_out);
    p9 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110101011010110101001101000100010011000100",
            TABLE => "0000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010010000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101100010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101101011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010011101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010011011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p9_in,
            y(0) => p9_out,
            y(1 to 14 - 1) => dummy9
        );


    p10_in <= x(8) & x(39) & x(59) & x(61) & x(62) & x(64) & x(65) & x(77) & x(90) & x(95) & x(101) & x(133) & x(149) & x(156) & x(164) & x(169) & x(171) & x(179) & x(200) & x(216) & x(227) & x(229) & x(233) & x(245) & x(251);
    y(10) <= not(p10_out);
    p10 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010010000110111110100100",
            TABLE => "0100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101101111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101101011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => 21,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p10_in,
            y(0) => p10_out,
            y(1 to 14 - 1) => dummy10
        );


    p11_in <= x(6) & x(10) & x(12) & x(23) & x(27) & x(34) & x(44) & x(46) & x(55) & x(61) & x(64) & x(73) & x(75) & x(79) & x(89) & x(101) & x(111) & x(118) & x(128) & x(132) & x(155) & x(156) & x(173) & x(177) & x(183) & x(194) & x(196) & x(206) & x(225) & x(242);
    y(11) <= not(p11_out);
    p11 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111011000011010101001110100110",
            TABLE => "000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 25,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p11_in,
            y(0) => p11_out,
            y(1 to 14 - 1) => dummy11
        );


    p12_in <= x(4) & x(5) & x(6) & x(27) & x(28) & x(35) & x(42) & x(46) & x(49) & x(51) & x(52) & x(53) & x(62) & x(72) & x(75) & x(77) & x(90) & x(103) & x(104) & x(111) & x(120) & x(130) & x(135) & x(143) & x(144) & x(149) & x(161) & x(172) & x(176) & x(177) & x(187) & x(194) & x(196) & x(210) & x(218) & x(231) & x(233) & x(236) & x(237) & x(245) & x(247) & x(248) & x(249) & x(251) & x(255);
    y(12) <= not(p12_out);
    p12 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110111000101111110111000110001110110010100010",
            TABLE => "000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001101100101001011011111111",
            SHIFT => 4,
            B => -47,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p12_in,
            y(0) => p12_out,
            y(1 to 15 - 1) => dummy12
        );


    p13_in <= x(4) & x(16) & x(21) & x(22) & x(29) & x(33) & x(38) & x(52) & x(53) & x(55) & x(60) & x(66) & x(69) & x(70) & x(103) & x(113) & x(133) & x(136) & x(137) & x(138) & x(141) & x(142) & x(143) & x(156) & x(161) & x(179) & x(180) & x(185) & x(188) & x(195) & x(222) & x(225) & x(230) & x(238) & x(244) & x(253);
    y(13) <= not(p13_out);
    p13 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101010100000000010100001000011011111",
            TABLE => "001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p13_in,
            y(0) => p13_out,
            y(1 to 15 - 1) => dummy13
        );


    p14_in <= x(1) & x(7) & x(18) & x(20) & x(22) & x(27) & x(30) & x(32) & x(33) & x(46) & x(65) & x(74) & x(89) & x(99) & x(100) & x(110) & x(127) & x(137) & x(142) & x(152) & x(154) & x(172) & x(173) & x(174) & x(176) & x(191) & x(204) & x(221) & x(225) & x(232) & x(236) & x(244) & x(245);
    y(14) <= not(p14_out);
    p14 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110001110010010001010110001110101",
            TABLE => "010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110010011010110100111111111",
            SHIFT => 4,
            B => 47,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p14_in,
            y(0) => p14_out,
            y(1 to 15 - 1) => dummy14
        );


    p15_in <= x(12) & x(16) & x(22) & x(30) & x(33) & x(35) & x(61) & x(65) & x(69) & x(74) & x(75) & x(78) & x(85) & x(93) & x(100) & x(106) & x(108) & x(111) & x(125) & x(127) & x(132) & x(134) & x(136) & x(149) & x(151) & x(152) & x(158) & x(166) & x(189) & x(213) & x(214) & x(225) & x(243);
    y(15) <= not(p15_out);
    p15 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000011110111111111111001100011011",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 4,
            B => -26,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p15_in,
            y(0) => p15_out,
            y(1 to 15 - 1) => dummy15
        );


    p16_in <= x(1) & x(7) & x(8) & x(12) & x(27) & x(34) & x(46) & x(50) & x(51) & x(55) & x(58) & x(62) & x(63) & x(75) & x(82) & x(89) & x(90) & x(119) & x(131) & x(133) & x(148) & x(151) & x(153) & x(167) & x(171) & x(177) & x(183) & x(189) & x(200) & x(213) & x(214) & x(218) & x(221) & x(229) & x(232) & x(250);
    y(16) <= not(p16_out);
    p16 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000110010000101110001000000000011",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 40,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p16_in,
            y(0) => p16_out,
            y(1 to 15 - 1) => dummy16
        );


    p17_in <= x(8) & x(14) & x(26) & x(33) & x(53) & x(55) & x(70) & x(111) & x(114) & x(120) & x(128) & x(139) & x(141) & x(158) & x(162) & x(165) & x(174) & x(175) & x(184) & x(201) & x(213) & x(221) & x(240) & x(242) & x(249) & x(255);
    y(17) <= not(p17_out);
    p17 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111111101111101001101101",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 4,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p17_in,
            y(0) => p17_out,
            y(1 to 14 - 1) => dummy17
        );


    p18_in <= x(6) & x(10) & x(18) & x(27) & x(33) & x(55) & x(61) & x(70) & x(76) & x(84) & x(93) & x(109) & x(111) & x(113) & x(118) & x(130) & x(143) & x(146) & x(156) & x(172) & x(181) & x(185) & x(187) & x(188) & x(195) & x(196) & x(204) & x(213) & x(225) & x(236) & x(238) & x(246);
    y(18) <= not(p18_out);
    p18 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101111101011001001111001010101",
            TABLE => "011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => -47,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p18_in,
            y(0) => p18_out,
            y(1 to 15 - 1) => dummy18
        );


    p19_in <= x(10) & x(16) & x(23) & x(39) & x(45) & x(52) & x(53) & x(77) & x(90) & x(106) & x(120) & x(127) & x(138) & x(139) & x(145) & x(147) & x(148) & x(156) & x(158) & x(165) & x(175) & x(181) & x(185) & x(190) & x(191) & x(219) & x(225) & x(226) & x(230) & x(234) & x(236) & x(241) & x(243) & x(244);
    y(19) <= not(p19_out);
    p19 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0101111010000110001001100001001010",
            TABLE => "0001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010011000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010011000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101101110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100010000010110010001001001011001001101001100101100000000000000000",
            SHIFT => 4,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p19_in,
            y(0) => p19_out,
            y(1 to 15 - 1) => dummy19
        );


    p20_in <= x(6) & x(29) & x(53) & x(61) & x(70) & x(78) & x(86) & x(109) & x(114) & x(126) & x(130) & x(147) & x(164) & x(168) & x(170) & x(171) & x(178) & x(181) & x(189) & x(191) & x(197) & x(201) & x(206) & x(208) & x(235) & x(236);
    y(20) <= not(p20_out);
    p20 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11010111101101110011111110",
            TABLE => "000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p20_in,
            y(0) => p20_out,
            y(1 to 14 - 1) => dummy20
        );


    p21_in <= x(4) & x(6) & x(10) & x(25) & x(58) & x(61) & x(62) & x(65) & x(70) & x(75) & x(89) & x(96) & x(98) & x(119) & x(131) & x(134) & x(136) & x(138) & x(149) & x(150) & x(155) & x(161) & x(174) & x(177) & x(178) & x(194) & x(197) & x(201) & x(223) & x(226) & x(231);
    y(21) <= not(p21_out);
    p21 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110110110110110110001101011011",
            TABLE => "0001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010011011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010010000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 25,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p21_in,
            y(0) => p21_out,
            y(1 to 15 - 1) => dummy21
        );


    p22_in <= x(2) & x(4) & x(21) & x(23) & x(27) & x(28) & x(29) & x(39) & x(41) & x(77) & x(79) & x(96) & x(99) & x(105) & x(112) & x(113) & x(114) & x(126) & x(129) & x(142) & x(143) & x(147) & x(149) & x(150) & x(162) & x(173) & x(203) & x(209) & x(229) & x(231) & x(238) & x(241) & x(243) & x(246) & x(248);
    y(22) <= not(p22_out);
    p22 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11110010110101001000011110110011011",
            TABLE => "00000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100100000100010011010000000000000100010011011101111100000100010011010010010001001101101100100010010001001101110110110010010001001101100101100110100101101001100101100110100110010110100101100110100110110010001000001111101110110010001000000000000010110010001000001011001000100100110110111011001000100100010011011011001000100100100101100110100101101001100101100110100110010110100101100110100101111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011000001000100011100000000000001000100011101110111100001000100011100001100010001110011100010001100010001110111001110001100010001110011010011001011010010110011010011001011001101001011010011001011000010000011100010111000111110111000110000111000101110001111001111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p22_in,
            y(0) => p22_out,
            y(1 to 15 - 1) => dummy22
        );


    p23_in <= x(5) & x(20) & x(30) & x(37) & x(47) & x(48) & x(77) & x(78) & x(81) & x(86) & x(88) & x(97) & x(100) & x(110) & x(112) & x(121) & x(122) & x(126) & x(135) & x(142) & x(147) & x(150) & x(160) & x(169) & x(170) & x(172) & x(188) & x(215) & x(216) & x(255);
    y(23) <= not(p23_out);
    p23 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110000100001111001010001001110",
            TABLE => "100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -48,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p23_in,
            y(0) => p23_out,
            y(1 to 14 - 1) => dummy23
        );


    p24_in <= x(0) & x(3) & x(23) & x(30) & x(38) & x(59) & x(66) & x(77) & x(78) & x(86) & x(96) & x(97) & x(98) & x(99) & x(100) & x(110) & x(112) & x(118) & x(127) & x(137) & x(143) & x(146) & x(148) & x(152) & x(164) & x(170) & x(172) & x(175) & x(177) & x(184) & x(195) & x(203) & x(204) & x(213) & x(215) & x(229) & x(237) & x(239) & x(252);
    y(24) <= not(p24_out);
    p24 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000101101100100001011011111101001001111",
            TABLE => "110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 4,
            B => 40,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p24_in,
            y(0) => p24_out,
            y(1 to 15 - 1) => dummy24
        );


    p25_in <= x(8) & x(10) & x(15) & x(29) & x(30) & x(31) & x(39) & x(42) & x(46) & x(51) & x(52) & x(54) & x(58) & x(65) & x(67) & x(79) & x(83) & x(88) & x(89) & x(91) & x(93) & x(115) & x(129) & x(138) & x(139) & x(144) & x(151) & x(161) & x(165) & x(166) & x(169) & x(170) & x(171) & x(173) & x(174) & x(184) & x(185) & x(198) & x(200) & x(201) & x(202) & x(206) & x(207) & x(211) & x(219) & x(220) & x(222) & x(225) & x(227) & x(234) & x(235) & x(242);
    y(25) <= not(p25_out);
    p25 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010010110110010111101001100011110100001111100100111",
            TABLE => "0100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101100000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101100100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101100000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101100001011100000001000101111000000110010110011010010000000000000000",
            SHIFT => 4,
            B => 19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p25_in,
            y(0) => p25_out,
            y(1 to 15 - 1) => dummy25
        );


    p26_in <= x(4) & x(17) & x(23) & x(36) & x(43) & x(47) & x(56) & x(72) & x(80) & x(97) & x(98) & x(100) & x(103) & x(119) & x(161) & x(168) & x(181) & x(194) & x(200) & x(211) & x(215) & x(223) & x(233) & x(239) & x(244);
    y(26) <= not(p26_out);
    p26 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100100001011111001010100",
            TABLE => "1011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010011101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010010000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => 52,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p26_in,
            y(0) => p26_out,
            y(1 to 14 - 1) => dummy26
        );


    p27_in <= x(0) & x(1) & x(7) & x(10) & x(23) & x(25) & x(38) & x(57) & x(91) & x(96) & x(105) & x(107) & x(117) & x(118) & x(119) & x(120) & x(125) & x(148) & x(150) & x(159) & x(161) & x(175) & x(179) & x(189) & x(212) & x(215) & x(233) & x(235) & x(238) & x(242) & x(250);
    y(27) <= not(p27_out);
    p27 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001101101101010000010001111111",
            TABLE => "1011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010010000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010011000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010011110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 33,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p27_in,
            y(0) => p27_out,
            y(1 to 15 - 1) => dummy27
        );


    p28_in <= x(6) & x(10) & x(14) & x(20) & x(25) & x(45) & x(55) & x(61) & x(96) & x(104) & x(105) & x(121) & x(126) & x(128) & x(129) & x(142) & x(152) & x(154) & x(158) & x(160) & x(163) & x(173) & x(188) & x(198) & x(208) & x(225) & x(226) & x(235) & x(244) & x(248) & x(252);
    y(28) <= not(p28_out);
    p28 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100000010110010100111001111001",
            TABLE => "1000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101101011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010010000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 63,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p28_in,
            y(0) => p28_out,
            y(1 to 15 - 1) => dummy28
        );


    p29_in <= x(15) & x(19) & x(35) & x(37) & x(41) & x(44) & x(47) & x(48) & x(51) & x(55) & x(61) & x(62) & x(75) & x(83) & x(95) & x(101) & x(112) & x(118) & x(121) & x(127) & x(143) & x(166) & x(169) & x(179) & x(194) & x(203) & x(216) & x(223) & x(229) & x(239) & x(242) & x(250) & x(255);
    y(29) <= not(p29_out);
    p29 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100011000000010110010110011000010",
            TABLE => "011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001101100101001011011111111",
            SHIFT => 4,
            B => 37,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p29_in,
            y(0) => p29_out,
            y(1 to 15 - 1) => dummy29
        );


    p30_in <= x(10) & x(27) & x(33) & x(46) & x(47) & x(55) & x(57) & x(70) & x(73) & x(83) & x(84) & x(98) & x(107) & x(109) & x(130) & x(137) & x(139) & x(152) & x(153) & x(156) & x(158) & x(168) & x(184) & x(188) & x(191) & x(193) & x(211) & x(213) & x(221) & x(222) & x(225) & x(230) & x(249);
    y(30) <= not(p30_out);
    p30 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001011010100000010101000001101000",
            TABLE => "011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 4,
            B => -36,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p30_in,
            y(0) => p30_out,
            y(1 to 15 - 1) => dummy30
        );


    p31_in <= x(4) & x(6) & x(8) & x(23) & x(44) & x(61) & x(63) & x(65) & x(68) & x(76) & x(78) & x(87) & x(93) & x(95) & x(96) & x(108) & x(114) & x(122) & x(125) & x(133) & x(139) & x(141) & x(143) & x(172) & x(178) & x(189) & x(195) & x(211) & x(226) & x(227) & x(235) & x(239) & x(243) & x(246) & x(247);
    y(31) <= not(p31_out);
    p31 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111010100101100000110000111010000",
            TABLE => "00000000000000100000001000101011000000100010101100101011101111111101010001000010010000100010101101000010001010110010101110111101011010011001011010010110011010011001011001101001011010011001011001000000110101000000000001000000110101001111110101000000110101000100001011010100001010110100001011010100101111010100001011010100011010011001011010010110011010011001011001101001011010011001011010000000111010001110100011111110000000001000000010000000111010001000000111101000111010000111111000010111100000011000000111101000100101100110100101101001100101100110100110010110100101100110100110001110111011110000100010001110000010001000111000000000000010001000111011100111000110001000111000011000100011100111000100011000100101100110100101101001100101100110100110010110100101100110100100101011101111110000001000101011000000100010101100000000000000100010101110111101010000100010101101000010001010111101010001000010011010011001011010010110011010011001011001101001011010011001011011101000100000001111111011101000111010001000000101111110111010000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 24,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p31_in,
            y(0) => p31_out,
            y(1 to 15 - 1) => dummy31
        );


    p32_in <= x(1) & x(2) & x(37) & x(48) & x(52) & x(56) & x(66) & x(75) & x(77) & x(93) & x(103) & x(110) & x(117) & x(120) & x(122) & x(134) & x(156) & x(167) & x(176) & x(179) & x(182) & x(187) & x(188) & x(189) & x(194) & x(215) & x(217) & x(238) & x(241) & x(243) & x(248) & x(251) & x(254);
    y(32) <= not(p32_out);
    p32 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101110110100001000010101101001000",
            TABLE => "000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p32_in,
            y(0) => p32_out,
            y(1 to 15 - 1) => dummy32
        );


    p33_in <= x(24) & x(30) & x(33) & x(36) & x(37) & x(46) & x(49) & x(55) & x(61) & x(72) & x(74) & x(102) & x(103) & x(105) & x(108) & x(114) & x(118) & x(127) & x(137) & x(142) & x(149) & x(157) & x(160) & x(173) & x(176) & x(178) & x(184) & x(188) & x(203) & x(215) & x(221) & x(226) & x(227) & x(228) & x(236) & x(241) & x(248) & x(250);
    y(33) <= not(p33_out);
    p33 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10101111101010100101100010011100010110",
            TABLE => "000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p33_in,
            y(0) => p33_out,
            y(1 to 15 - 1) => dummy33
        );


    p34_in <= x(5) & x(10) & x(14) & x(23) & x(25) & x(31) & x(32) & x(34) & x(45) & x(47) & x(49) & x(54) & x(55) & x(64) & x(70) & x(77) & x(83) & x(109) & x(116) & x(118) & x(122) & x(123) & x(128) & x(133) & x(135) & x(139) & x(143) & x(165) & x(171) & x(172) & x(185) & x(191) & x(195) & x(196) & x(200) & x(202) & x(218) & x(221) & x(234) & x(238) & x(241) & x(243) & x(250) & x(251) & x(252) & x(255);
    y(34) <= not(p34_out);
    p34 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101010000000101111001011001101110111111101100",
            TABLE => "0000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010010100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100000100010001110000110001000111001101001100101100000000000000000",
            SHIFT => 4,
            B => -17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p34_in,
            y(0) => p34_out,
            y(1 to 15 - 1) => dummy34
        );


    p35_in <= x(3) & x(25) & x(30) & x(36) & x(43) & x(55) & x(56) & x(73) & x(89) & x(91) & x(97) & x(134) & x(154) & x(159) & x(161) & x(171) & x(173) & x(174) & x(193) & x(194) & x(196) & x(199) & x(200) & x(215) & x(219) & x(226) & x(231) & x(234) & x(244) & x(248);
    y(35) <= not(p35_out);
    p35 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000110111101010101110100000110",
            TABLE => "101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 5,
            B => -24,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p35_in,
            y(0) => p35_out,
            y(1 to 15 - 1) => dummy35
        );


    p36_in <= x(1) & x(4) & x(10) & x(31) & x(47) & x(68) & x(69) & x(75) & x(77) & x(91) & x(96) & x(106) & x(108) & x(127) & x(148) & x(149) & x(150) & x(156) & x(157) & x(161) & x(162) & x(177) & x(189) & x(194) & x(198) & x(209) & x(226) & x(229) & x(231) & x(233) & x(250);
    y(36) <= not(p36_out);
    p36 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0011011000100000001110000011111",
            TABLE => "0100110111011111000001000100110100000100010011010000000000000100010011011101101100100100010011010010010001001101101100100010010001101001100101101001011001101001100101100110100101101001100101101011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 24,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p36_in,
            y(0) => p36_out,
            y(1 to 15 - 1) => dummy36
        );


    p37_in <= x(13) & x(15) & x(27) & x(35) & x(39) & x(40) & x(41) & x(48) & x(53) & x(57) & x(61) & x(62) & x(80) & x(89) & x(95) & x(107) & x(109) & x(110) & x(118) & x(125) & x(127) & x(128) & x(129) & x(138) & x(139) & x(158) & x(166) & x(169) & x(172) & x(177) & x(188) & x(197) & x(202) & x(216) & x(219) & x(231) & x(254) & x(255);
    y(37) <= not(p37_out);
    p37 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10111101011101100011011100001101001111",
            TABLE => "000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 4,
            B => -28,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p37_in,
            y(0) => p37_out,
            y(1 to 15 - 1) => dummy37
        );


    p38_in <= x(4) & x(6) & x(10) & x(13) & x(25) & x(36) & x(37) & x(40) & x(47) & x(53) & x(55) & x(56) & x(65) & x(69) & x(71) & x(73) & x(77) & x(78) & x(80) & x(83) & x(89) & x(91) & x(93) & x(100) & x(105) & x(106) & x(142) & x(143) & x(156) & x(158) & x(172) & x(179) & x(180) & x(190) & x(193) & x(195) & x(196) & x(200) & x(225) & x(238) & x(244) & x(248);
    y(38) <= not(p38_out);
    p38 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000011111111011001101100001101111010100011",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p38_in,
            y(0) => p38_out,
            y(1 to 15 - 1) => dummy38
        );


    p39_in <= x(8) & x(10) & x(22) & x(27) & x(31) & x(32) & x(33) & x(44) & x(61) & x(64) & x(68) & x(74) & x(83) & x(89) & x(98) & x(109) & x(112) & x(116) & x(120) & x(124) & x(139) & x(162) & x(165) & x(173) & x(174) & x(177) & x(184) & x(189) & x(201) & x(202) & x(211) & x(220) & x(221) & x(222) & x(225) & x(226) & x(227) & x(236) & x(239) & x(251);
    y(39) <= not(p39_out);
    p39 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010101110111100100011001101111001010000",
            TABLE => "0010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101100000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101101000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101101110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p39_in,
            y(0) => p39_out,
            y(1 to 15 - 1) => dummy39
        );


    p40_in <= x(8) & x(17) & x(20) & x(21) & x(25) & x(30) & x(35) & x(42) & x(44) & x(49) & x(57) & x(61) & x(64) & x(89) & x(95) & x(100) & x(101) & x(116) & x(117) & x(121) & x(126) & x(133) & x(137) & x(142) & x(154) & x(174) & x(179) & x(182) & x(191) & x(204) & x(208) & x(209) & x(225) & x(226) & x(244) & x(255);
    y(40) <= not(p40_out);
    p40 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001110001111110111101101110110010010",
            TABLE => "001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -49,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p40_in,
            y(0) => p40_out,
            y(1 to 15 - 1) => dummy40
        );


    p41_in <= x(26) & x(38) & x(52) & x(53) & x(69) & x(76) & x(121) & x(145) & x(148) & x(155) & x(156) & x(166) & x(183) & x(185) & x(189) & x(194) & x(196) & x(202) & x(203) & x(210) & x(224) & x(227) & x(246) & x(255);
    y(41) <= not(p41_out);
    p41 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000101000000011111110110",
            TABLE => "110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p41_in,
            y(0) => p41_out,
            y(1 to 14 - 1) => dummy41
        );


    p42_in <= x(22) & x(30) & x(40) & x(52) & x(61) & x(65) & x(83) & x(89) & x(93) & x(100) & x(102) & x(128) & x(129) & x(130) & x(137) & x(138) & x(159) & x(160) & x(161) & x(165) & x(173) & x(174) & x(176) & x(184) & x(221) & x(225) & x(236) & x(238) & x(244) & x(250);
    y(42) <= not(p42_out);
    p42 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100110110101010010000110000010",
            TABLE => "001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -55,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p42_in,
            y(0) => p42_out,
            y(1 to 15 - 1) => dummy42
        );


    p43_in <= x(7) & x(11) & x(21) & x(23) & x(24) & x(26) & x(33) & x(38) & x(40) & x(49) & x(61) & x(71) & x(72) & x(79) & x(88) & x(89) & x(102) & x(103) & x(111) & x(120) & x(136) & x(142) & x(144) & x(157) & x(161) & x(173) & x(175) & x(198) & x(201) & x(210) & x(212) & x(215) & x(220) & x(225) & x(231) & x(233) & x(249);
    y(43) <= not(p43_out);
    p43 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010110011010100010111001111000111111",
            TABLE => "0001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010010100110111011111000001000100110100000100010011010000000000000100010011011101101100100100010011010010010001001101101100100010010001101001100101101001011001101001100101100110100101101001100101101101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010010000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p43_in,
            y(0) => p43_out,
            y(1 to 15 - 1) => dummy43
        );


    p44_in <= x(7) & x(11) & x(22) & x(23) & x(30) & x(33) & x(40) & x(44) & x(61) & x(64) & x(77) & x(80) & x(81) & x(83) & x(89) & x(92) & x(97) & x(100) & x(101) & x(110) & x(119) & x(137) & x(149) & x(152) & x(154) & x(168) & x(173) & x(176) & x(179) & x(189) & x(212) & x(221) & x(225) & x(227) & x(244) & x(252);
    y(44) <= not(p44_out);
    p44 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100010100101100000100101001010011011",
            TABLE => "101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 43,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p44_in,
            y(0) => p44_out,
            y(1 to 15 - 1) => dummy44
        );


    p45_in <= x(5) & x(21) & x(31) & x(38) & x(39) & x(41) & x(46) & x(48) & x(60) & x(66) & x(88) & x(96) & x(97) & x(102) & x(112) & x(118) & x(140) & x(170) & x(172) & x(179) & x(196) & x(215) & x(222) & x(226) & x(235) & x(237) & x(240) & x(245) & x(246) & x(247);
    y(45) <= not(p45_out);
    p45 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110011010001101010000100000111",
            TABLE => "000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -52,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p45_in,
            y(0) => p45_out,
            y(1 to 14 - 1) => dummy45
        );


    p46_in <= x(2) & x(3) & x(6) & x(8) & x(12) & x(33) & x(38) & x(62) & x(76) & x(77) & x(78) & x(91) & x(104) & x(121) & x(139) & x(149) & x(167) & x(171) & x(182) & x(187) & x(189) & x(196) & x(232) & x(233) & x(247);
    y(46) <= not(p46_out);
    p46 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000010111110101001111000",
            TABLE => "1111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101101000111000001000111011111000111000001000000000001000111000001000100011100001100011100111100011100001100001110001100011100001100010010110011010010110100110010110011010011001011010010110011010010000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -49,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p46_in,
            y(0) => p46_out,
            y(1 to 14 - 1) => dummy46
        );


    p47_in <= x(1) & x(2) & x(7) & x(16) & x(27) & x(30) & x(43) & x(50) & x(52) & x(54) & x(68) & x(70) & x(72) & x(75) & x(81) & x(91) & x(96) & x(99) & x(106) & x(108) & x(112) & x(113) & x(122) & x(125) & x(130) & x(139) & x(149) & x(165) & x(167) & x(174) & x(179) & x(189) & x(194) & x(196) & x(200) & x(218) & x(223) & x(226) & x(233) & x(239);
    y(47) <= not(p47_out);
    p47 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010111011000111011100110011001111111001",
            TABLE => "0001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010010000100010001110000000000000100010001110111011110000100010001110000110001000111001110001000110001000111011100111000110001000111001101001100101101001011001101001100101100110100101101001100101100000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010011000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010100000011010100010000101101010001101001100101100000000000000000",
            SHIFT => 4,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p47_in,
            y(0) => p47_out,
            y(1 to 15 - 1) => dummy47
        );


    p48_in <= x(3) & x(10) & x(28) & x(29) & x(35) & x(53) & x(61) & x(62) & x(71) & x(78) & x(80) & x(105) & x(113) & x(126) & x(128) & x(130) & x(135) & x(147) & x(148) & x(156) & x(169) & x(179) & x(189) & x(191) & x(196) & x(213) & x(214) & x(225) & x(229) & x(236) & x(254);
    y(48) <= not(p48_out);
    p48 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001001011010011110001111000100",
            TABLE => "1110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101101011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p48_in,
            y(0) => p48_out,
            y(1 to 15 - 1) => dummy48
        );


    p49_in <= x(6) & x(10) & x(14) & x(25) & x(27) & x(29) & x(33) & x(39) & x(44) & x(46) & x(53) & x(55) & x(61) & x(70) & x(75) & x(81) & x(97) & x(111) & x(131) & x(135) & x(137) & x(142) & x(147) & x(152) & x(156) & x(163) & x(165) & x(173) & x(177) & x(180) & x(181) & x(184) & x(185) & x(194) & x(195) & x(213) & x(225) & x(237) & x(243) & x(248) & x(253);
    y(49) <= not(p49_out);
    p49 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00110011101111101100010000001110110100110",
            TABLE => "10001110111011110000100010001110000010001000111000000000000010001000111011100111000110001000111000011000100011100111000100011000100101100110100101101001100101100110100110010110100101100110100100000000000100000001000001110001000100000111000101110001111101111000111000011000000110000111000100011000011100010111000111100111011010011001011010010110011010011001011001101001011010011001011000000000000100000001000001110001000100000111000101110001111101111000111000011000000110000111000100011000011100010111000111100111011010011001011010010110011010011001011001101001011010011001011011101111100011101000111000001000100011100000100000001000000000001110011110001110100011100001100010001110000110000001100001110001011010011001011010010110011010011001011001101001011010011001011011110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100100000100010011010000000000000100010011011101111100000100010011010010010001001101101100100010010001001101110110110010010001001101100101100110100101101001100101100110100110010110100101100110100110111111001010110010101100000010101111010010101100101011010000101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -67,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p49_in,
            y(0) => p49_out,
            y(1 to 15 - 1) => dummy49
        );


    p50_in <= x(4) & x(8) & x(13) & x(18) & x(29) & x(57) & x(83) & x(84) & x(85) & x(94) & x(95) & x(103) & x(107) & x(109) & x(129) & x(139) & x(140) & x(141) & x(142) & x(154) & x(168) & x(178) & x(189) & x(191) & x(203) & x(211) & x(222) & x(226) & x(228) & x(230) & x(235) & x(244) & x(247) & x(254);
    y(50) <= not(p50_out);
    p50 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111001010100011110000100111101001",
            TABLE => "0000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010010100000011010100010000101101010001101001100101100000000000000000",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p50_in,
            y(0) => p50_out,
            y(1 to 15 - 1) => dummy50
        );


    p51_in <= x(7) & x(11) & x(12) & x(14) & x(17) & x(18) & x(39) & x(45) & x(50) & x(66) & x(76) & x(77) & x(78) & x(80) & x(88) & x(95) & x(99) & x(106) & x(111) & x(118) & x(146) & x(152) & x(174) & x(177) & x(195) & x(196) & x(208) & x(218) & x(225) & x(235) & x(236) & x(238) & x(241) & x(250) & x(251);
    y(51) <= not(p51_out);
    p51 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10101000000100011100110110111101101",
            TABLE => "00100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011011111101110101001101010001000000110101000100000001000000000000001011110111010100110101000100001011010100010000100100001000101011011010011001011010010110011010011001011001101001011010011001011001111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011001001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011000000001000101110000000000000001000101110111111100000001000101111000000100010111111010001000000100010111011111101000000100010111011010011001011010010110011010011001011001101001011010011001011001001101110111110000010001001101010011011101101100100100010011010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p51_in,
            y(0) => p51_out,
            y(1 to 15 - 1) => dummy51
        );


    p52_in <= x(10) & x(27) & x(44) & x(46) & x(61) & x(72) & x(80) & x(82) & x(91) & x(95) & x(99) & x(100) & x(114) & x(142) & x(158) & x(161) & x(179) & x(187) & x(215) & x(231) & x(248);
    y(52) <= not(p52_out);
    p52 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110110000111010110111",
            TABLE => "000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => 4,
            B => 16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p52_in,
            y(0) => p52_out,
            y(1 to 14 - 1) => dummy52
        );


    p53_in <= x(7) & x(8) & x(10) & x(13) & x(24) & x(25) & x(30) & x(43) & x(53) & x(61) & x(66) & x(67) & x(79) & x(88) & x(105) & x(117) & x(119) & x(120) & x(148) & x(156) & x(158) & x(162) & x(171) & x(174) & x(192) & x(193) & x(195) & x(198) & x(201) & x(203) & x(220) & x(225) & x(236) & x(242) & x(250);
    y(53) <= not(p53_out);
    p53 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10111110000010000111000000110011000",
            TABLE => "00000001000101110000000000000001000101110111111100000001000101111000000100010111111010001000000100010111011111101000000100010111011010011001011010010110011010011001011001101001011010011001011011101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011011010100010000000100000000000000111111011101010011010100010000001101010001000010010000100010101110111101110101001101010001000010100101100110100101101001100101100110100110010110100101100110100110000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100110001110111011110000100010001110000010001000111000000000000010001000111011100111000110001000111000011000100011100111000100011000100101100110100101101001100101100110100110010110100101100110100110000000111010001110100011111110100000011110100011101000011111101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -27,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p53_in,
            y(0) => p53_out,
            y(1 to 15 - 1) => dummy53
        );


    p54_in <= x(4) & x(10) & x(16) & x(17) & x(23) & x(25) & x(27) & x(29) & x(32) & x(33) & x(34) & x(38) & x(78) & x(90) & x(93) & x(97) & x(102) & x(112) & x(136) & x(138) & x(142) & x(143) & x(156) & x(157) & x(158) & x(171) & x(180) & x(181) & x(214) & x(215) & x(217) & x(225) & x(230) & x(234) & x(239) & x(248) & x(250) & x(253);
    y(54) <= not(p54_out);
    p54 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11001011000110101001001101000001110011",
            TABLE => "001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 4,
            B => 29,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p54_in,
            y(0) => p54_out,
            y(1 to 15 - 1) => dummy54
        );


    p55_in <= x(1) & x(21) & x(22) & x(23) & x(30) & x(44) & x(48) & x(57) & x(61) & x(77) & x(92) & x(97) & x(100) & x(110) & x(119) & x(121) & x(125) & x(137) & x(142) & x(154) & x(155) & x(158) & x(168) & x(172) & x(173) & x(177) & x(191) & x(203) & x(215) & x(218) & x(241) & x(248) & x(252) & x(255);
    y(55) <= not(p55_out);
    p55 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000101000000001010001011000000011",
            TABLE => "1011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010011101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101100111000100010000011100010001100001101001100101100000000000000000",
            SHIFT => 4,
            B => 50,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p55_in,
            y(0) => p55_out,
            y(1 to 15 - 1) => dummy55
        );


    p56_in <= x(1) & x(5) & x(6) & x(10) & x(57) & x(63) & x(64) & x(68) & x(77) & x(84) & x(87) & x(89) & x(93) & x(95) & x(96) & x(100) & x(101) & x(102) & x(104) & x(115) & x(134) & x(140) & x(146) & x(150) & x(164) & x(169) & x(189) & x(192) & x(199) & x(225) & x(226) & x(228) & x(231) & x(235) & x(238) & x(241) & x(247);
    y(56) <= not(p56_out);
    p56 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100001000001000111001011111110100001",
            TABLE => "1000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101100111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101100100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 3,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p56_in,
            y(0) => p56_out,
            y(1 to 14 - 1) => dummy56
        );


    p57_in <= x(2) & x(7) & x(13) & x(28) & x(29) & x(35) & x(39) & x(54) & x(61) & x(66) & x(78) & x(80) & x(88) & x(91) & x(96) & x(112) & x(116) & x(119) & x(128) & x(130) & x(159) & x(163) & x(167) & x(170) & x(179) & x(181) & x(185) & x(188) & x(190) & x(201) & x(212) & x(217) & x(225) & x(227) & x(230) & x(234) & x(244) & x(250) & x(255);
    y(57) <= not(p57_out);
    p57 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000111101000001011100110011000110100110",
            TABLE => "011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110001010110110100111111111",
            SHIFT => 4,
            B => -20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p57_in,
            y(0) => p57_out,
            y(1 to 15 - 1) => dummy57
        );


    p58_in <= x(1) & x(4) & x(23) & x(33) & x(45) & x(48) & x(58) & x(67) & x(78) & x(92) & x(99) & x(101) & x(114) & x(119) & x(128) & x(132) & x(143) & x(146) & x(155) & x(156) & x(161) & x(166) & x(173) & x(177) & x(178) & x(183) & x(185) & x(191) & x(195) & x(206) & x(211) & x(222) & x(228) & x(236) & x(241);
    y(58) <= not(p58_out);
    p58 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001010100111111000101010100000010",
            TABLE => "11111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011001000000110101000000000001000000110101001111110101000000110101000100001011010100001010110100001011010100101111010100001011010100011010011001011010010110011010011001011001101001011010011001011000000000000000100000001000101011000000100010101100101011101111111101010001000010010000100010101101000010001010110010101110111101011010011001011010010110011010011001011001101001011010011001011010110010111110110010000010110010001000001011001000000000001000001011001011011011001001001011001000100100101100100100110100100100100101100110100101101001100101100110100110010110100101100110100110000000111010000000000010000000111010001111111010000000111010001000000111101000000101111000000111101000011111101000000111101000100101100110100101101001100101100110100110010110100101100110100111111011101100101011001000100000110110111011001010110010001001000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p58_in,
            y(0) => p58_out,
            y(1 to 15 - 1) => dummy58
        );


    p59_in <= x(6) & x(7) & x(27) & x(30) & x(33) & x(34) & x(41) & x(51) & x(52) & x(54) & x(65) & x(92) & x(94) & x(95) & x(106) & x(110) & x(112) & x(114) & x(142) & x(166) & x(169) & x(197) & x(207) & x(229) & x(238) & x(248) & x(250);
    y(59) <= not(p59_out);
    p59 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000010101101100110111010001",
            TABLE => "111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001110101001001011011111111",
            SHIFT => 4,
            B => -28,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p59_in,
            y(0) => p59_out,
            y(1 to 14 - 1) => dummy59
        );


    p60_in <= x(10) & x(28) & x(35) & x(40) & x(41) & x(46) & x(57) & x(62) & x(65) & x(84) & x(101) & x(113) & x(121) & x(130) & x(132) & x(139) & x(155) & x(166) & x(173) & x(174) & x(178) & x(180) & x(182) & x(216) & x(217) & x(218) & x(226) & x(227) & x(231) & x(243) & x(248) & x(254);
    y(60) <= not(p60_out);
    p60 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001100001001011101000100000000",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => 19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p60_in,
            y(0) => p60_out,
            y(1 to 15 - 1) => dummy60
        );


    p61_in <= x(25) & x(61) & x(66) & x(69) & x(78) & x(85) & x(97) & x(98) & x(100) & x(126) & x(130) & x(143) & x(152) & x(154) & x(159) & x(160) & x(166) & x(169) & x(171) & x(176) & x(177) & x(183) & x(186) & x(189) & x(191) & x(208) & x(210) & x(216) & x(225) & x(235) & x(236) & x(241) & x(244) & x(246) & x(248) & x(250) & x(253);
    y(61) <= not(p61_out);
    p61 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101101010110110100111111100000111100",
            TABLE => "0000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010010001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010010010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101101000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -54,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p61_in,
            y(0) => p61_out,
            y(1 to 15 - 1) => dummy61
        );


    p62_in <= x(4) & x(5) & x(6) & x(25) & x(29) & x(31) & x(42) & x(43) & x(57) & x(61) & x(64) & x(84) & x(89) & x(91) & x(95) & x(111) & x(114) & x(115) & x(127) & x(140) & x(148) & x(155) & x(159) & x(162) & x(169) & x(170) & x(189) & x(208) & x(212) & x(226) & x(229) & x(231) & x(233) & x(235) & x(237) & x(238) & x(240) & x(253);
    y(62) <= not(p62_out);
    p62 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101111110110101100000101011111111110",
            TABLE => "011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => 40,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p62_in,
            y(0) => p62_out,
            y(1 to 15 - 1) => dummy62
        );


    p63_in <= x(6) & x(13) & x(25) & x(38) & x(43) & x(46) & x(53) & x(61) & x(73) & x(82) & x(89) & x(103) & x(107) & x(109) & x(114) & x(117) & x(119) & x(156) & x(167) & x(168) & x(169) & x(177) & x(179) & x(188) & x(189) & x(191) & x(194) & x(203) & x(211) & x(215) & x(216) & x(222) & x(229) & x(242) & x(250) & x(253);
    y(63) <= not(p63_out);
    p63 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111100010010000001000110101010011100",
            TABLE => "000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p63_in,
            y(0) => p63_out,
            y(1 to 15 - 1) => dummy63
        );


    p64_in <= x(1) & x(28) & x(35) & x(39) & x(44) & x(46) & x(52) & x(53) & x(69) & x(72) & x(77) & x(78) & x(93) & x(99) & x(102) & x(103) & x(107) & x(108) & x(129) & x(132) & x(142) & x(149) & x(164) & x(168) & x(169) & x(175) & x(176) & x(181) & x(191) & x(194) & x(202) & x(220) & x(226) & x(237) & x(244) & x(249) & x(254);
    y(64) <= not(p64_out);
    p64 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111100101101110001101000001011010001",
            TABLE => "0000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101101101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010011000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p64_in,
            y(0) => p64_out,
            y(1 to 15 - 1) => dummy64
        );


    p65_in <= x(2) & x(27) & x(34) & x(38) & x(46) & x(48) & x(58) & x(59) & x(91) & x(99) & x(103) & x(109) & x(117) & x(138) & x(139) & x(154) & x(156) & x(171) & x(174) & x(183) & x(189) & x(203) & x(210) & x(215) & x(227) & x(240) & x(247);
    y(65) <= not(p65_out);
    p65 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101001000010110000011101111",
            TABLE => "010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 5,
            B => -32,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p65_in,
            y(0) => p65_out,
            y(1 to 15 - 1) => dummy65
        );


    p66_in <= x(10) & x(25) & x(30) & x(34) & x(35) & x(55) & x(78) & x(80) & x(91) & x(95) & x(96) & x(97) & x(100) & x(109) & x(134) & x(138) & x(141) & x(148) & x(151) & x(159) & x(162) & x(164) & x(191) & x(194) & x(203) & x(226) & x(239) & x(243) & x(253);
    y(66) <= not(p66_out);
    p66 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10011100011110011010100011010",
            TABLE => "00010111000000010000000100000000011111110001011100010111000000010001011110000001100000011110100001111110000101110001011110000001100101100110100101101001100101100110100110010110100101100110100101111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011000101011000000100000001000000000101111110010101100101011000000100010101101000010010000101101010010111101001010110010101101000010011010011001011010010110011010011001011001101001011010011001011010000000111010000000000010000000111010001111111010000000111010001000000111101000000101111000000111101000011111101000000111101000100101100110100101101001100101100110100110010110100101100110100100100000101100101011001011111011001001001011001010110010110110110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 42,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p66_in,
            y(0) => p66_out,
            y(1 to 14 - 1) => dummy66
        );


    p67_in <= x(7) & x(10) & x(11) & x(18) & x(30) & x(33) & x(40) & x(61) & x(64) & x(80) & x(89) & x(92) & x(100) & x(101) & x(103) & x(117) & x(119) & x(120) & x(121) & x(128) & x(129) & x(136) & x(137) & x(148) & x(149) & x(156) & x(160) & x(162) & x(167) & x(168) & x(173) & x(177) & x(179) & x(184) & x(197) & x(203) & x(212) & x(220) & x(225) & x(241) & x(248);
    y(67) <= not(p67_out);
    p67 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00110101001110111001000010011101001110011",
            TABLE => "01001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011001110001000100001111011101110001000100000000000001110001000100000111000100011000111001110111000100011000100011100111000100011000011010011001011010010110011010011001011001101001011010011001011000000010001010110000000000000010001010111011111100000010001010110100001000101011110101000100001000101011101111010100001000101011100101100110100101101001100101100110100110010110100101100110100111101000100000001111111011101000100000000000000011101000100000001110100010000001011111101110100010000001000101111110100010000001011010011001011010010110011010011001011001101001011010011001011000010111000000010000000100000000011111110001011100010111000000010001011110000001100000011110100001111110000101110001011110000001100101100110100101101001100101100110100110010110100101100110100101110001000100001111011101110001000100000000000001110001000100000111000100011000111001110111000100011000100011100111000100011000011010011001011010010110011010011001011001101001011010011001011001110001000100001111011101110001011100010001100011100111011100010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p67_in,
            y(0) => p67_out,
            y(1 to 15 - 1) => dummy67
        );


    p68_in <= x(6) & x(7) & x(12) & x(14) & x(17) & x(33) & x(40) & x(61) & x(71) & x(76) & x(78) & x(96) & x(111) & x(116) & x(117) & x(119) & x(126) & x(128) & x(136) & x(143) & x(158) & x(162) & x(185) & x(195) & x(196) & x(199) & x(203) & x(209) & x(225) & x(231) & x(235) & x(236) & x(239) & x(243) & x(244) & x(249);
    y(68) <= not(p68_out);
    p68 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000101010110111111011110111100011110",
            TABLE => "110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -36,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p68_in,
            y(0) => p68_out,
            y(1 to 15 - 1) => dummy68
        );


    p69_in <= x(3) & x(10) & x(35) & x(38) & x(39) & x(46) & x(55) & x(72) & x(78) & x(80) & x(81) & x(87) & x(90) & x(91) & x(94) & x(96) & x(97) & x(99) & x(104) & x(114) & x(129) & x(135) & x(138) & x(143) & x(156) & x(170) & x(181) & x(193) & x(195) & x(196) & x(206) & x(226) & x(229) & x(249);
    y(69) <= not(p69_out);
    p69 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111100100011001111010101010100100",
            TABLE => "0000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101100010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101101000111000001000100011100001100010010110011010010000000000000000",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p69_in,
            y(0) => p69_out,
            y(1 to 15 - 1) => dummy69
        );


    p70_in <= x(6) & x(9) & x(12) & x(20) & x(28) & x(30) & x(35) & x(38) & x(45) & x(58) & x(65) & x(71) & x(76) & x(81) & x(96) & x(97) & x(100) & x(112) & x(114) & x(130) & x(138) & x(139) & x(157) & x(158) & x(165) & x(171) & x(172) & x(174) & x(176) & x(184) & x(196) & x(217) & x(225) & x(227) & x(233) & x(236) & x(249) & x(254);
    y(70) <= not(p70_out);
    p70 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001110111011000010101110100111110101",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => -28,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p70_in,
            y(0) => p70_out,
            y(1 to 15 - 1) => dummy70
        );


    p71_in <= x(9) & x(25) & x(27) & x(44) & x(45) & x(53) & x(56) & x(61) & x(65) & x(66) & x(67) & x(72) & x(154) & x(156) & x(161) & x(166) & x(171) & x(178) & x(179) & x(180) & x(182) & x(196) & x(199) & x(203) & x(204) & x(210) & x(220) & x(231) & x(233) & x(240) & x(248) & x(252);
    y(71) <= not(p71_out);
    p71 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01011001100010100101110100111110",
            TABLE => "001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => -29,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p71_in,
            y(0) => p71_out,
            y(1 to 15 - 1) => dummy71
        );


    p72_in <= x(6) & x(19) & x(27) & x(38) & x(44) & x(46) & x(54) & x(55) & x(56) & x(76) & x(81) & x(91) & x(96) & x(99) & x(103) & x(117) & x(122) & x(161) & x(179) & x(193) & x(199) & x(212) & x(220) & x(221) & x(223) & x(226) & x(231) & x(233) & x(238);
    y(72) <= not(p72_out);
    p72 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10001000000010110100011001111",
            TABLE => "10110010001000000010000000000000111110111011001010110010001000001011001000100100001001000100110111011011101100101011001000100100100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100000100010011010000000000000100010011011101111100000100010011010010010001001101101100100010010001001101110110110010010001001101100101100110100101101001100101100110100110010110100101100110100110111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100100010111011111110000000100010111000101110111111010000001000101111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p72_in,
            y(0) => p72_out,
            y(1 to 14 - 1) => dummy72
        );


    p73_in <= x(18) & x(37) & x(38) & x(44) & x(50) & x(70) & x(78) & x(81) & x(82) & x(87) & x(88) & x(89) & x(93) & x(98) & x(100) & x(102) & x(107) & x(109) & x(112) & x(114) & x(121) & x(127) & x(132) & x(137) & x(143) & x(152) & x(156) & x(203) & x(212) & x(221) & x(226) & x(229) & x(232);
    y(73) <= not(p73_out);
    p73 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010000111000010011011001110001010",
            TABLE => "111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => 4,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p73_in,
            y(0) => p73_out,
            y(1 to 15 - 1) => dummy73
        );


    p74_in <= x(27) & x(29) & x(42) & x(55) & x(69) & x(84) & x(95) & x(109) & x(111) & x(117) & x(132) & x(141) & x(142) & x(148) & x(156) & x(171) & x(174) & x(189) & x(191) & x(194) & x(200) & x(201) & x(202) & x(228) & x(244) & x(248) & x(250);
    y(74) <= not(p74_out);
    p74 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011011010100100110100110111",
            TABLE => "000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p74_in,
            y(0) => p74_out,
            y(1 to 14 - 1) => dummy74
        );


    p75_in <= x(0) & x(6) & x(7) & x(37) & x(39) & x(47) & x(62) & x(63) & x(73) & x(93) & x(95) & x(101) & x(105) & x(108) & x(112) & x(114) & x(121) & x(122) & x(124) & x(127) & x(129) & x(134) & x(142) & x(144) & x(156) & x(166) & x(167) & x(169) & x(172) & x(177) & x(194) & x(209) & x(214) & x(216) & x(230) & x(231) & x(248) & x(250) & x(253) & x(255);
    y(75) <= not(p75_out);
    p75 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000000011011110000100100111000001100110",
            TABLE => "1110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101100100110111011111000001000100110100000100010011010000000000000100010011011101101100100100010011010010010001001101101100100010010001101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101101011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010010000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101101011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010010010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p75_in,
            y(0) => p75_out,
            y(1 to 15 - 1) => dummy75
        );


    p76_in <= x(7) & x(10) & x(11) & x(13) & x(21) & x(34) & x(35) & x(65) & x(80) & x(82) & x(89) & x(90) & x(93) & x(95) & x(99) & x(124) & x(125) & x(127) & x(151) & x(154) & x(161) & x(168) & x(174) & x(176) & x(177) & x(183) & x(188) & x(197) & x(204) & x(214) & x(215) & x(229) & x(235) & x(242) & x(245);
    y(76) <= not(p76_out);
    p76 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101000101010000101001100000000000",
            TABLE => "10110010111110110010000010110010001000001011001000000000001000001011001011011011001001001011001000100100101100100100110100100100100101100110100101101001100101100110100110010110100101100110100110110010111110110010000010110010001000001011001000000000001000001011001011011011001001001011001000100100101100100100110100100100100101100110100101101001100101100110100110010110100101100110100111010100010000000100000000000000111111011101010011010100010000001101010001000010010000100010101110111101110101001101010001000010100101100110100101101001100101100110100110010110100101100110100101110001000100001111011101110001000100000000000001110001000100000111000100011000111001110111000100011000100011100111000100011000011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p76_in,
            y(0) => p76_out,
            y(1 to 15 - 1) => dummy76
        );


    p77_in <= x(13) & x(29) & x(55) & x(77) & x(88) & x(91) & x(95) & x(109) & x(111) & x(112) & x(147) & x(169) & x(172) & x(186) & x(191) & x(192) & x(195) & x(199) & x(209) & x(213) & x(218) & x(228) & x(230) & x(238) & x(241) & x(248);
    y(77) <= not(p77_out);
    p77 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10101100110110010101011000",
            TABLE => "000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p77_in,
            y(0) => p77_out,
            y(1 to 14 - 1) => dummy77
        );


    p78_in <= x(3) & x(31) & x(34) & x(35) & x(50) & x(56) & x(70) & x(75) & x(90) & x(107) & x(119) & x(127) & x(133) & x(135) & x(147) & x(151) & x(154) & x(156) & x(177) & x(189) & x(191) & x(192) & x(198) & x(214) & x(226) & x(227) & x(230) & x(232) & x(236) & x(242) & x(243) & x(244) & x(245);
    y(78) <= not(p78_out);
    p78 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101100111000000100110101110011101",
            TABLE => "000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001010011010110100111111111",
            SHIFT => 4,
            B => -27,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p78_in,
            y(0) => p78_out,
            y(1 to 15 - 1) => dummy78
        );


    p79_in <= x(17) & x(30) & x(36) & x(38) & x(45) & x(52) & x(56) & x(70) & x(97) & x(102) & x(103) & x(110) & x(118) & x(142) & x(156) & x(169) & x(176) & x(181) & x(183) & x(194) & x(203) & x(233);
    y(79) <= not(p79_out);
    p79 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111101001001010010100",
            TABLE => "0000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010011000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101101000111000001000100011100001100010010110011010010000000000000000",
            SHIFT => 5,
            B => 27,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p79_in,
            y(0) => p79_out,
            y(1 to 15 - 1) => dummy79
        );


    p80_in <= x(9) & x(16) & x(22) & x(25) & x(27) & x(29) & x(30) & x(65) & x(71) & x(73) & x(75) & x(78) & x(79) & x(93) & x(98) & x(105) & x(112) & x(113) & x(117) & x(130) & x(134) & x(136) & x(137) & x(142) & x(143) & x(144) & x(155) & x(162) & x(176) & x(207) & x(210) & x(221) & x(225) & x(229) & x(236) & x(238) & x(244) & x(248);
    y(80) <= not(p80_out);
    p80 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11110000100010001101110110101100000011",
            TABLE => "000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 4,
            B => -34,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p80_in,
            y(0) => p80_out,
            y(1 to 15 - 1) => dummy80
        );


    p81_in <= x(1) & x(4) & x(10) & x(27) & x(37) & x(45) & x(49) & x(52) & x(53) & x(68) & x(71) & x(80) & x(82) & x(87) & x(91) & x(93) & x(100) & x(111) & x(129) & x(143) & x(149) & x(150) & x(169) & x(172) & x(175) & x(179) & x(181) & x(189) & x(191) & x(193) & x(194) & x(196) & x(200) & x(206) & x(221) & x(226) & x(235) & x(236) & x(238) & x(242) & x(244) & x(249);
    y(81) <= not(p81_out);
    p81 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101110110011101001010111110111010110000011",
            TABLE => "000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p81_in,
            y(0) => p81_out,
            y(1 to 15 - 1) => dummy81
        );


    p82_in <= x(31) & x(39) & x(40) & x(43) & x(53) & x(54) & x(57) & x(61) & x(65) & x(77) & x(83) & x(117) & x(122) & x(127) & x(137) & x(148) & x(156) & x(162) & x(168) & x(174) & x(176) & x(185) & x(189) & x(203) & x(218) & x(221) & x(225) & x(227) & x(229) & x(232) & x(236) & x(248);
    y(82) <= not(p82_out);
    p82 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000100001011011001100000100100",
            TABLE => "111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => 22,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p82_in,
            y(0) => p82_out,
            y(1 to 15 - 1) => dummy82
        );


    p83_in <= x(2) & x(5) & x(24) & x(27) & x(30) & x(34) & x(35) & x(55) & x(58) & x(61) & x(66) & x(93) & x(96) & x(101) & x(118) & x(121) & x(139) & x(143) & x(146) & x(164) & x(169) & x(170) & x(174) & x(176) & x(193) & x(203) & x(206) & x(215) & x(229) & x(233) & x(239) & x(255);
    y(83) <= not(p83_out);
    p83 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11100000000111001011101101010100",
            TABLE => "000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p83_in,
            y(0) => p83_out,
            y(1 to 15 - 1) => dummy83
        );


    p84_in <= x(7) & x(14) & x(16) & x(17) & x(36) & x(39) & x(46) & x(48) & x(52) & x(56) & x(64) & x(70) & x(72) & x(73) & x(85) & x(98) & x(103) & x(111) & x(117) & x(130) & x(134) & x(141) & x(145) & x(146) & x(156) & x(166) & x(168) & x(169) & x(183) & x(207) & x(213) & x(215) & x(221) & x(239) & x(246);
    y(84) <= not(p84_out);
    p84 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10110010100001001001111111111111000",
            TABLE => "00001000100011100000000000001000100011101110111100001000100011100001100010001110011100010001100010001110111001110001100010001110011010011001011010010110011010011001011001101001011010011001011010000000111010000000000010000000111010001111111010000000111010001000000111101000000101111000000111101000011111101000000111101000100101100110100101101001100101100110100110010110100101100110100110110010001000001111101110110010001000000000000010110010001000001011001000100100110110111011001000100100010011011011001000100100100101100110100101101001100101100110100110010110100101100110100100000001000101110001011101111111000000000000000100000001000101111000000100010111000101110111111011101000100000011000000100010111011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100110000000111010001110100011111110100000011110100011101000011111101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p84_in,
            y(0) => p84_out,
            y(1 to 15 - 1) => dummy84
        );


    p85_in <= x(2) & x(5) & x(13) & x(41) & x(53) & x(55) & x(61) & x(73) & x(77) & x(83) & x(109) & x(117) & x(119) & x(145) & x(152) & x(156) & x(169) & x(188) & x(196) & x(199) & x(200) & x(203) & x(211) & x(216) & x(222) & x(229);
    y(85) <= not(p85_out);
    p85 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00100110010001010010001011",
            TABLE => "110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 4,
            B => -20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p85_in,
            y(0) => p85_out,
            y(1 to 14 - 1) => dummy85
        );


    p86_in <= x(0) & x(12) & x(17) & x(22) & x(24) & x(29) & x(36) & x(46) & x(48) & x(53) & x(56) & x(59) & x(61) & x(62) & x(69) & x(79) & x(86) & x(89) & x(93) & x(97) & x(98) & x(102) & x(105) & x(110) & x(112) & x(114) & x(117) & x(121) & x(127) & x(135) & x(137) & x(153) & x(155) & x(156) & x(161) & x(169) & x(171) & x(178) & x(194) & x(200) & x(212) & x(215) & x(221) & x(228) & x(229) & x(233) & x(244) & x(250);
    y(86) <= not(p86_out);
    p86 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000001101111111011001110011101100000111010101011",
            TABLE => "111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p86_in,
            y(0) => p86_out,
            y(1 to 15 - 1) => dummy86
        );


    p87_in <= x(6) & x(8) & x(10) & x(14) & x(18) & x(22) & x(23) & x(33) & x(45) & x(53) & x(55) & x(57) & x(70) & x(77) & x(88) & x(97) & x(103) & x(112) & x(114) & x(120) & x(126) & x(128) & x(131) & x(137) & x(141) & x(142) & x(156) & x(158) & x(159) & x(160) & x(169) & x(176) & x(184) & x(191) & x(195) & x(197) & x(198) & x(199) & x(203) & x(207) & x(221) & x(225) & x(231) & x(236) & x(238) & x(242) & x(244) & x(247);
    y(87) <= not(p87_out);
    p87 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010111011110101111001100110100110000011100010101",
            TABLE => "000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p87_in,
            y(0) => p87_out,
            y(1 to 15 - 1) => dummy87
        );


    p88_in <= x(7) & x(10) & x(11) & x(18) & x(19) & x(25) & x(33) & x(35) & x(49) & x(50) & x(70) & x(87) & x(89) & x(91) & x(99) & x(102) & x(137) & x(138) & x(142) & x(152) & x(155) & x(156) & x(159) & x(194) & x(226) & x(234) & x(253);
    y(88) <= not(p88_out);
    p88 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011110110111100101000110110",
            TABLE => "000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001001010110110100111111111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p88_in,
            y(0) => p88_out,
            y(1 to 14 - 1) => dummy88
        );


    p89_in <= x(18) & x(26) & x(27) & x(35) & x(37) & x(39) & x(45) & x(46) & x(49) & x(60) & x(61) & x(70) & x(80) & x(85) & x(91) & x(92) & x(94) & x(109) & x(111) & x(117) & x(130) & x(132) & x(146) & x(147) & x(148) & x(155) & x(156) & x(159) & x(166) & x(185) & x(187) & x(204) & x(213) & x(220) & x(227) & x(236) & x(242) & x(243) & x(246) & x(247);
    y(89) <= not(p89_out);
    p89 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001011010110100001101000000011011111111",
            TABLE => "0100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010011110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101100000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101101111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 4,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p89_in,
            y(0) => p89_out,
            y(1 to 15 - 1) => dummy89
        );


    p90_in <= x(2) & x(5) & x(26) & x(27) & x(44) & x(55) & x(59) & x(60) & x(76) & x(83) & x(91) & x(96) & x(114) & x(137) & x(141) & x(150) & x(156) & x(171) & x(178) & x(196) & x(201) & x(202) & x(239);
    y(90) <= not(p90_out);
    p90 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11101000010101000110110",
            TABLE => "00000000001000000010000010110010001000001011001010110010111110110100110100100100001001001011001000100100101100101011001011011011100101100110100101101001100101100110100110010110100101100110100111011111010011010100110100000100010011010000010000000100000000001101101101001101010011010010010001001101001001000010010010110010100101100110100101101001100101100110100110010110100101100110100111010100010000001111110111010100010000000000000011010100010000001101010001000010101111011101010001000010001010111101010001000010100101100110100101101001100101100110100110010110100101100110100100101011000000101011111100101011001010110100001010111101001010110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 5,
            B => 17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p90_in,
            y(0) => p90_out,
            y(1 to 15 - 1) => dummy90
        );


    p91_in <= x(8) & x(10) & x(17) & x(18) & x(22) & x(26) & x(36) & x(39) & x(49) & x(56) & x(59) & x(81) & x(92) & x(98) & x(99) & x(102) & x(104) & x(114) & x(120) & x(143) & x(148) & x(149) & x(154) & x(156) & x(166) & x(172) & x(175) & x(180) & x(189) & x(203) & x(213) & x(215) & x(234) & x(235) & x(247) & x(249) & x(253);
    y(91) <= not(p91_out);
    p91 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010110000001011101000101001010111000",
            TABLE => "0001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010011011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010010100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p91_in,
            y(0) => p91_out,
            y(1 to 15 - 1) => dummy91
        );


    p92_in <= x(6) & x(7) & x(8) & x(13) & x(24) & x(33) & x(35) & x(47) & x(49) & x(72) & x(88) & x(89) & x(101) & x(102) & x(111) & x(120) & x(142) & x(161) & x(173) & x(192) & x(200) & x(215) & x(217) & x(220) & x(231) & x(247) & x(249);
    y(92) <= not(p92_out);
    p92 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001001110111011000010000000",
            TABLE => "110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 4,
            B => -33,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p92_in,
            y(0) => p92_out,
            y(1 to 14 - 1) => dummy92
        );


    p93_in <= x(10) & x(25) & x(29) & x(47) & x(48) & x(65) & x(72) & x(85) & x(91) & x(111) & x(113) & x(132) & x(139) & x(140) & x(159) & x(161) & x(168) & x(194) & x(200) & x(230) & x(233) & x(238) & x(248);
    y(93) <= not(p93_out);
    p93 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10100100001000011010111",
            TABLE => "01000000110101000000000001000000110101001111110101000000110101000100001011010100001010110100001011010100101111010100001011010100011010011001011010010110011010011001011001101001011010011001011011111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011010111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100100010111000000010111111100010111000101111000000101111110000101111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 51,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p93_in,
            y(0) => p93_out,
            y(1 to 14 - 1) => dummy93
        );


    p94_in <= x(8) & x(14) & x(19) & x(28) & x(37) & x(56) & x(70) & x(97) & x(113) & x(135) & x(137) & x(142) & x(143) & x(147) & x(156) & x(164) & x(170) & x(189) & x(194) & x(205) & x(213) & x(215) & x(229) & x(237) & x(241) & x(243) & x(248);
    y(94) <= not(p94_out);
    p94 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011101111001101100011100011",
            TABLE => "000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 4,
            B => -31,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p94_in,
            y(0) => p94_out,
            y(1 to 14 - 1) => dummy94
        );


    p95_in <= x(6) & x(13) & x(27) & x(33) & x(34) & x(45) & x(47) & x(55) & x(61) & x(64) & x(70) & x(72) & x(89) & x(93) & x(99) & x(121) & x(137) & x(138) & x(152) & x(154) & x(163) & x(167) & x(171) & x(180) & x(183) & x(186) & x(195) & x(202) & x(204) & x(214) & x(219) & x(221) & x(225) & x(229) & x(240) & x(248) & x(249) & x(250) & x(253) & x(255);
    y(95) <= not(p95_out);
    p95 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000000001010100101011100011100110001110",
            TABLE => "1110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010011011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010010000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010010101110111111000000100010101100000010001010110000000000000010001010111011110101000010001010110100001000101011110101000100001001101001100101101001011001101001100101100110100101101001100101101000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010000001000101011010000100010101110010110011010010000000000000000",
            SHIFT => 4,
            B => 30,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p95_in,
            y(0) => p95_out,
            y(1 to 15 - 1) => dummy95
        );


    p96_in <= x(1) & x(10) & x(23) & x(25) & x(35) & x(36) & x(38) & x(42) & x(78) & x(80) & x(87) & x(91) & x(95) & x(100) & x(107) & x(110) & x(120) & x(138) & x(143) & x(145) & x(155) & x(167) & x(171) & x(191) & x(198) & x(223) & x(226) & x(235) & x(239) & x(242) & x(249);
    y(96) <= not(p96_out);
    p96 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001010011010010101010011100101",
            TABLE => "0100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100100110111011111000001000100110100000100010011010000000000000100010011011101101100100100010011010010010001001101101100100010010001101001100101101001011001101001100101100110100101101001100101101011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010010100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => -48,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p96_in,
            y(0) => p96_out,
            y(1 to 15 - 1) => dummy96
        );


    p97_in <= x(4) & x(10) & x(23) & x(27) & x(34) & x(39) & x(41) & x(114) & x(124) & x(127) & x(138) & x(143) & x(149) & x(161) & x(173) & x(177) & x(178) & x(184) & x(202) & x(203) & x(211) & x(217) & x(222) & x(225) & x(227) & x(231) & x(236);
    y(97) <= not(p97_out);
    p97 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101000100100100100101010000",
            TABLE => "100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 4,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p97_in,
            y(0) => p97_out,
            y(1 to 14 - 1) => dummy97
        );


    p98_in <= x(47) & x(56) & x(61) & x(62) & x(76) & x(77) & x(79) & x(81) & x(84) & x(96) & x(114) & x(156) & x(161) & x(169) & x(187) & x(215) & x(226) & x(231) & x(233) & x(239) & x(244) & x(253);
    y(98) <= not(p98_out);
    p98 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111110110110010000110",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010011110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 5,
            B => -43,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p98_in,
            y(0) => p98_out,
            y(1 to 15 - 1) => dummy98
        );


    p99_in <= x(23) & x(27) & x(44) & x(52) & x(60) & x(66) & x(73) & x(75) & x(95) & x(96) & x(97) & x(98) & x(100) & x(110) & x(112) & x(122) & x(128) & x(137) & x(146) & x(156) & x(164) & x(171) & x(177) & x(182) & x(185) & x(199) & x(202) & x(203) & x(211) & x(215) & x(222) & x(233) & x(235) & x(236) & x(254);
    y(99) <= not(p99_out);
    p99 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10101000111011100011001100011111101",
            TABLE => "00100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011000101011101111110000001000101011000000100010101100000000000000100010101110111101010000100010101101000010001010111101010001000010011010011001011010010110011010011001011001101001011010011001011000000000100000001000000011101000100000001110100011101000111111100001011110000001100000011110100010000001111010001110100001111110011010011001011010010110011010011001011001101001011010011001011000010000000000000111000100010000011100010001000011110111011100010001100010001110011100010001100001110001000110001110011101110001100101100110100101101001100101100110100110010110100101100110100101111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011000000100010011010100110111011111001001000100110101001101110110111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -38,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p99_in,
            y(0) => p99_out,
            y(1 to 15 - 1) => dummy99
        );


    p100_in <= x(3) & x(17) & x(31) & x(32) & x(34) & x(37) & x(49) & x(59) & x(93) & x(109) & x(113) & x(122) & x(127) & x(143) & x(163) & x(164) & x(177) & x(180) & x(183) & x(191) & x(210) & x(213) & x(214) & x(224) & x(235) & x(243) & x(250) & x(253);
    y(100) <= not(p100_out);
    p100 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010000111001011000110000011",
            TABLE => "1110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000100010001110000000000000100010001110111011110000100010001110000110001000111001110001000110001000111011100111000110001000111001101001100101101001011001101001100101100110100101101001100101101000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010111000100010000011100010001100001101001100101100000000000000000",
            SHIFT => 4,
            B => 37,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p100_in,
            y(0) => p100_out,
            y(1 to 14 - 1) => dummy100
        );


    p101_in <= x(3) & x(6) & x(7) & x(17) & x(21) & x(22) & x(31) & x(37) & x(40) & x(43) & x(50) & x(53) & x(71) & x(76) & x(95) & x(98) & x(99) & x(137) & x(143) & x(153) & x(155) & x(157) & x(158) & x(167) & x(174) & x(177) & x(183) & x(185) & x(191) & x(193) & x(196) & x(199) & x(212) & x(214) & x(215) & x(218) & x(222) & x(228) & x(236) & x(244) & x(248) & x(250);
    y(101) <= not(p101_out);
    p101 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111101011000101010011000011000000111110010",
            TABLE => "000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p101_in,
            y(0) => p101_out,
            y(1 to 15 - 1) => dummy101
        );


    p102_in <= x(5) & x(30) & x(33) & x(50) & x(54) & x(56) & x(61) & x(70) & x(77) & x(93) & x(109) & x(121) & x(141) & x(150) & x(155) & x(167) & x(172) & x(175) & x(179) & x(187) & x(188) & x(189) & x(196) & x(211) & x(214) & x(222) & x(238) & x(241);
    y(102) <= not(p102_out);
    p102 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001010010100001000010000011",
            TABLE => "0100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101101011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010011110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101101110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100111000100010000011100010001100001101001100101100000000000000000",
            SHIFT => 4,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p102_in,
            y(0) => p102_out,
            y(1 to 14 - 1) => dummy102
        );


    p103_in <= x(4) & x(5) & x(10) & x(13) & x(18) & x(20) & x(27) & x(31) & x(34) & x(35) & x(42) & x(55) & x(58) & x(65) & x(69) & x(77) & x(82) & x(111) & x(115) & x(118) & x(121) & x(124) & x(127) & x(135) & x(161) & x(168) & x(169) & x(173) & x(174) & x(177) & x(184) & x(202) & x(208) & x(213) & x(221) & x(225) & x(226) & x(236) & x(241);
    y(103) <= not(p103_out);
    p103 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001100111111111000111101110100101011110",
            TABLE => "100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001001010110110100111111111",
            SHIFT => 4,
            B => 22,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p103_in,
            y(0) => p103_out,
            y(1 to 15 - 1) => dummy103
        );


    p104_in <= x(4) & x(29) & x(32) & x(33) & x(36) & x(37) & x(55) & x(61) & x(65) & x(67) & x(74) & x(87) & x(91) & x(105) & x(114) & x(117) & x(127) & x(134) & x(136) & x(156) & x(158) & x(162) & x(172) & x(179) & x(193) & x(195) & x(196) & x(201) & x(203) & x(204) & x(212) & x(239) & x(241) & x(246);
    y(104) <= not(p104_out);
    p104 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100000110110111100001000101101011",
            TABLE => "1000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010011110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101100001000001110001000110000111000110010110011010010000000000000000",
            SHIFT => 4,
            B => -20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p104_in,
            y(0) => p104_out,
            y(1 to 15 - 1) => dummy104
        );


    p105_in <= x(5) & x(10) & x(29) & x(30) & x(54) & x(59) & x(72) & x(75) & x(86) & x(99) & x(109) & x(111) & x(114) & x(127) & x(132) & x(143) & x(147) & x(156) & x(161) & x(168) & x(177) & x(179) & x(185) & x(189) & x(194) & x(195) & x(203) & x(206) & x(208) & x(225) & x(231) & x(244);
    y(105) <= not(p105_out);
    p105 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01111100101011011111010001011111",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 4,
            B => 15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p105_in,
            y(0) => p105_out,
            y(1 to 15 - 1) => dummy105
        );


    p106_in <= x(13) & x(23) & x(24) & x(29) & x(42) & x(43) & x(61) & x(62) & x(77) & x(78) & x(79) & x(80) & x(86) & x(87) & x(89) & x(92) & x(105) & x(107) & x(109) & x(113) & x(117) & x(126) & x(135) & x(136) & x(142) & x(145) & x(147) & x(156) & x(168) & x(173) & x(189) & x(191) & x(197) & x(213) & x(225) & x(236) & x(254);
    y(106) <= not(p106_out);
    p106 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101111111001011111010100011101110000",
            TABLE => "0000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101100010101110111111000000100010101100000010001010110000000000000010001010111011110101000010001010110100001000101011110101000100001001101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p106_in,
            y(0) => p106_out,
            y(1 to 15 - 1) => dummy106
        );


    p107_in <= x(2) & x(6) & x(7) & x(23) & x(31) & x(44) & x(45) & x(50) & x(52) & x(56) & x(57) & x(58) & x(71) & x(76) & x(80) & x(83) & x(86) & x(88) & x(95) & x(96) & x(117) & x(152) & x(166) & x(185) & x(187) & x(188) & x(191) & x(193) & x(200) & x(204) & x(220) & x(225) & x(233) & x(235) & x(239) & x(246) & x(247) & x(251);
    y(107) <= not(p107_out);
    p107 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00011101111101111100101110110000001100",
            TABLE => "011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => -53,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p107_in,
            y(0) => p107_out,
            y(1 to 15 - 1) => dummy107
        );


    p108_in <= x(0) & x(2) & x(3) & x(20) & x(25) & x(38) & x(39) & x(49) & x(55) & x(62) & x(72) & x(75) & x(77) & x(81) & x(91) & x(93) & x(95) & x(97) & x(101) & x(110) & x(112) & x(114) & x(120) & x(129) & x(141) & x(142) & x(165) & x(176) & x(180) & x(187) & x(208) & x(226) & x(228) & x(235) & x(242) & x(247) & x(248);
    y(108) <= not(p108_out);
    p108 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000001001111101100101010010011101100",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010010100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101101101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010010000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => 28,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p108_in,
            y(0) => p108_out,
            y(1 to 15 - 1) => dummy108
        );


    p109_in <= x(19) & x(29) & x(32) & x(44) & x(48) & x(53) & x(62) & x(76) & x(78) & x(90) & x(108) & x(121) & x(124) & x(127) & x(136) & x(156) & x(158) & x(176) & x(181) & x(185) & x(190) & x(201) & x(233) & x(236);
    y(109) <= not(p109_out);
    p109 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010110001010010101001110",
            TABLE => "001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p109_in,
            y(0) => p109_out,
            y(1 to 15 - 1) => dummy109
        );


    p110_in <= x(2) & x(4) & x(25) & x(33) & x(38) & x(43) & x(49) & x(53) & x(61) & x(62) & x(80) & x(96) & x(103) & x(111) & x(115) & x(142) & x(148) & x(150) & x(151) & x(156) & x(157) & x(158) & x(161) & x(162) & x(168) & x(195) & x(198) & x(203) & x(213) & x(225) & x(230) & x(232) & x(235) & x(238) & x(240) & x(242) & x(244) & x(248) & x(254) & x(255);
    y(110) <= not(p110_out);
    p110 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110101000100100111100000110111100001000",
            TABLE => "0010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101101011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010010111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101101000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010011000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011000000011101000100000011110100010010110011010010000000000000000",
            SHIFT => 4,
            B => -49,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p110_in,
            y(0) => p110_out,
            y(1 to 15 - 1) => dummy110
        );


    p111_in <= x(23) & x(24) & x(32) & x(34) & x(37) & x(43) & x(45) & x(49) & x(55) & x(74) & x(76) & x(77) & x(97) & x(99) & x(104) & x(107) & x(119) & x(123) & x(127) & x(130) & x(133) & x(135) & x(165) & x(166) & x(172) & x(180) & x(186) & x(187) & x(189) & x(191) & x(210) & x(231) & x(234) & x(238) & x(247) & x(250);
    y(111) <= not(p111_out);
    p111 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100001000111000111101111001101101101",
            TABLE => "110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p111_in,
            y(0) => p111_out,
            y(1 to 15 - 1) => dummy111
        );


    p112_in <= x(27) & x(35) & x(48) & x(52) & x(58) & x(72) & x(87) & x(89) & x(93) & x(103) & x(108) & x(127) & x(129) & x(137) & x(139) & x(140) & x(142) & x(144) & x(154) & x(156) & x(168) & x(171) & x(176) & x(191) & x(194) & x(198) & x(203) & x(210) & x(215) & x(221) & x(232) & x(235) & x(241) & x(242) & x(244) & x(248);
    y(112) <= not(p112_out);
    p112 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111001101000111101010100100101110100",
            TABLE => "000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 23,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p112_in,
            y(0) => p112_out,
            y(1 to 15 - 1) => dummy112
        );


    p113_in <= x(1) & x(4) & x(8) & x(17) & x(24) & x(36) & x(45) & x(46) & x(61) & x(72) & x(83) & x(103) & x(108) & x(111) & x(113) & x(114) & x(124) & x(126) & x(138) & x(139) & x(140) & x(141) & x(142) & x(150) & x(154) & x(161) & x(168) & x(169) & x(177) & x(178) & x(187) & x(188) & x(193) & x(194) & x(203) & x(211) & x(212) & x(215) & x(216) & x(220) & x(225) & x(232);
    y(113) <= not(p113_out);
    p113 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111001001110010000011101000010100101000001",
            TABLE => "000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p113_in,
            y(0) => p113_out,
            y(1 to 15 - 1) => dummy113
        );


    p114_in <= x(10) & x(11) & x(27) & x(32) & x(33) & x(44) & x(52) & x(56) & x(60) & x(61) & x(62) & x(65) & x(70) & x(82) & x(98) & x(104) & x(114) & x(122) & x(142) & x(152) & x(154) & x(165) & x(174) & x(176) & x(199) & x(201) & x(204) & x(211) & x(222) & x(225) & x(232) & x(236) & x(244) & x(246) & x(252);
    y(114) <= not(p114_out);
    p114 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01001111110010000010101101011010110",
            TABLE => "01110001000100001111011101110001000100000000000001110001000100000111000100011000111001110111000100011000100011100111000100011000011010011001011010010110011010011001011001101001011010011001011000000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100111101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011000010000011100010000000000010000011100011111011100010000011100010001100001110001100011100001100001110001111001110001100001110001100101100110100101101001100101100110100110010110100101100110100100101011000000101011111100101011000000100000000000101011000000100010101101000010101111010010101101000010110101000010101101000010011010011001011010010110011010011001011001101001011010011001011000101011000000101011111100101011001010110100001010111101001010110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -57,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p114_in,
            y(0) => p114_out,
            y(1 to 15 - 1) => dummy114
        );


    p115_in <= x(2) & x(4) & x(8) & x(10) & x(56) & x(62) & x(72) & x(76) & x(78) & x(87) & x(91) & x(93) & x(113) & x(139) & x(141) & x(156) & x(158) & x(173) & x(185) & x(190) & x(196) & x(213) & x(215) & x(220) & x(225) & x(226) & x(251);
    y(115) <= not(p115_out);
    p115 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111100100101011100010001111",
            TABLE => "000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 4,
            B => 21,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p115_in,
            y(0) => p115_out,
            y(1 to 14 - 1) => dummy115
        );


    p116_in <= x(5) & x(10) & x(35) & x(38) & x(45) & x(46) & x(47) & x(53) & x(54) & x(76) & x(78) & x(86) & x(99) & x(111) & x(114) & x(124) & x(126) & x(128) & x(139) & x(141) & x(147) & x(153) & x(156) & x(164) & x(165) & x(166) & x(171) & x(176) & x(184) & x(185) & x(195) & x(207) & x(233) & x(234) & x(236) & x(253);
    y(116) <= not(p116_out);
    p116 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110100000000110011110111001100101001",
            TABLE => "000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p116_in,
            y(0) => p116_out,
            y(1 to 15 - 1) => dummy116
        );


    p117_in <= x(17) & x(19) & x(22) & x(27) & x(38) & x(43) & x(46) & x(59) & x(61) & x(79) & x(81) & x(97) & x(110) & x(112) & x(121) & x(122) & x(130) & x(138) & x(155) & x(158) & x(169) & x(179) & x(196) & x(203) & x(233) & x(239);
    y(117) <= not(p117_out);
    p117 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01011111101000110101011001",
            TABLE => "000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => 28,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p117_in,
            y(0) => p117_out,
            y(1 to 14 - 1) => dummy117
        );


    p118_in <= x(1) & x(3) & x(7) & x(11) & x(12) & x(14) & x(16) & x(27) & x(41) & x(62) & x(68) & x(73) & x(87) & x(88) & x(89) & x(90) & x(98) & x(120) & x(125) & x(128) & x(156) & x(174) & x(175) & x(186) & x(189) & x(197) & x(200) & x(201) & x(218) & x(223) & x(226) & x(227) & x(232) & x(233) & x(245);
    y(118) <= not(p118_out);
    p118 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11101001110100011110001110101101001",
            TABLE => "00000000001000000010000010110010001000001011001010110010111110110100110100100100001001001011001000100100101100101011001011011011100101100110100101101001100101100110100110010110100101100110100100000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100101111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011001110001000100000001000000000000111101110111000101110001000100000111000100011000000110001000111011100111011100010111000100011000011010011001011010010110011010011001011001101001011010011001011000010000011100010000000000010000011100011111011100010000011100010001100001110001100011100001100001110001111001110001100001110001100101100110100101101001100101100110100110010110100101100110100111010100111111010100000011010100110101001011110101000010110101001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p118_in,
            y(0) => p118_out,
            y(1 to 15 - 1) => dummy118
        );


    p119_in <= x(6) & x(10) & x(17) & x(18) & x(22) & x(34) & x(48) & x(64) & x(68) & x(70) & x(75) & x(76) & x(78) & x(81) & x(89) & x(96) & x(97) & x(98) & x(125) & x(149) & x(176) & x(182) & x(189) & x(201) & x(203) & x(212) & x(223) & x(226) & x(233) & x(239);
    y(119) <= not(p119_out);
    p119 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111011001100001110001101110110",
            TABLE => "000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p119_in,
            y(0) => p119_out,
            y(1 to 14 - 1) => dummy119
        );


    p120_in <= x(1) & x(10) & x(14) & x(24) & x(27) & x(31) & x(32) & x(39) & x(65) & x(70) & x(88) & x(103) & x(107) & x(109) & x(111) & x(122) & x(124) & x(132) & x(135) & x(137) & x(139) & x(147) & x(156) & x(157) & x(191) & x(192) & x(206) & x(221) & x(230) & x(249);
    y(120) <= not(p120_out);
    p120 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110011001010110010110111101101",
            TABLE => "000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p120_in,
            y(0) => p120_out,
            y(1 to 14 - 1) => dummy120
        );


    p121_in <= x(2) & x(25) & x(35) & x(48) & x(52) & x(53) & x(64) & x(68) & x(69) & x(70) & x(77) & x(85) & x(90) & x(109) & x(111) & x(115) & x(130) & x(138) & x(166) & x(168) & x(171) & x(176) & x(183) & x(193) & x(202) & x(225);
    y(121) <= not(p121_out);
    p121 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11010010010100100100010001",
            TABLE => "000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p121_in,
            y(0) => p121_out,
            y(1 to 14 - 1) => dummy121
        );


    p122_in <= x(6) & x(8) & x(11) & x(12) & x(24) & x(47) & x(53) & x(54) & x(72) & x(79) & x(83) & x(88) & x(100) & x(120) & x(130) & x(139) & x(158) & x(161) & x(187) & x(200) & x(242) & x(249);
    y(122) <= not(p122_out);
    p122 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001100001001110010101",
            TABLE => "0010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101101110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010010100110100000100010011010010010001101001100101100000000000000000",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p122_in,
            y(0) => p122_out,
            y(1 to 15 - 1) => dummy122
        );


    p123_in <= x(0) & x(12) & x(22) & x(26) & x(28) & x(30) & x(46) & x(48) & x(65) & x(68) & x(100) & x(110) & x(112) & x(114) & x(121) & x(130) & x(137) & x(142) & x(169) & x(173) & x(174) & x(176) & x(185) & x(188) & x(215) & x(228) & x(229) & x(236) & x(239);
    y(123) <= not(p123_out);
    p123 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001101100001101001001000111",
            TABLE => "11110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100110000000111010001110100011111110000000001000000010000000111010001000000111101000111010000111111000010111100000011000000111101000100101100110100101101001100101100110100110010110100101100110100100100000101100101011001011111011000000000010000000100000101100100010010010110010101100101101101101001101001001000010010010110010011010011001011010010110011010011001011001101001011010011001011010110010001000001111101110110010001000000000000010110010001000001011001000100100110110111011001000100100010011011011001000100100100101100110100101101001100101100110100110010110100101100110100101111111000101110001011100000001011111100001011100010111100000010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p123_in,
            y(0) => p123_out,
            y(1 to 14 - 1) => dummy123
        );


    p124_in <= x(6) & x(13) & x(22) & x(24) & x(33) & x(44) & x(46) & x(47) & x(52) & x(56) & x(91) & x(94) & x(95) & x(96) & x(127) & x(129) & x(131) & x(132) & x(145) & x(151) & x(154) & x(160) & x(161) & x(168) & x(169) & x(173) & x(189) & x(221) & x(223) & x(224) & x(235) & x(238);
    y(124) <= not(p124_out);
    p124 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00111011101100100000100110000100",
            TABLE => "001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p124_in,
            y(0) => p124_out,
            y(1 to 15 - 1) => dummy124
        );


    p125_in <= x(4) & x(20) & x(52) & x(56) & x(61) & x(69) & x(77) & x(90) & x(91) & x(105) & x(113) & x(142) & x(143) & x(172) & x(179) & x(181) & x(187) & x(193) & x(195) & x(221) & x(225) & x(226) & x(234) & x(238) & x(239);
    y(125) <= not(p125_out);
    p125 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000001101000001101011110",
            TABLE => "1110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101100000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101101011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010010000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p125_in,
            y(0) => p125_out,
            y(1 to 14 - 1) => dummy125
        );


    p126_in <= x(4) & x(5) & x(7) & x(10) & x(13) & x(23) & x(32) & x(34) & x(40) & x(44) & x(55) & x(77) & x(82) & x(83) & x(109) & x(121) & x(122) & x(127) & x(132) & x(137) & x(143) & x(150) & x(172) & x(175) & x(179) & x(195) & x(196) & x(202) & x(204) & x(219) & x(230) & x(250) & x(251) & x(255);
    y(126) <= not(p126_out);
    p126 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100010001011110011000000101001110",
            TABLE => "0100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101101101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010010000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101000111000001000111011111000111000001000000000001000111000001000100011100001100011100111100011100001100001110001100011100001100010010110011010010110100110010110011010011001011010010110011010010000001000101011010000100010101110010110011010010000000000000000",
            SHIFT => 4,
            B => -34,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p126_in,
            y(0) => p126_out,
            y(1 to 15 - 1) => dummy126
        );


    p127_in <= x(12) & x(13) & x(23) & x(29) & x(37) & x(45) & x(52) & x(54) & x(65) & x(70) & x(85) & x(89) & x(90) & x(92) & x(101) & x(115) & x(118) & x(128) & x(134) & x(135) & x(150) & x(168) & x(174) & x(191) & x(218) & x(225) & x(236) & x(244) & x(254);
    y(127) <= not(p127_out);
    p127 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10111010000101010111111110010",
            TABLE => "00000010001010110000000000000010001010111011111100000010001010110100001000101011110101000100001000101011101111010100001000101011100101100110100101101001100101100110100110010110100101100110100111010100010000000100000000000000111111011101010011010100010000001101010001000010010000100010101110111101110101001101010001000010100101100110100101101001100101100110100110010110100101100110100101001101000001001101111101001101000001000000000001001101000001000100110100100100110110110100110100100100101100100100110100100100011010011001011010010110011010011001011001101001011010011001011000000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100110110010001000001111101110110010101100100010010011011011101100101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p127_in,
            y(0) => p127_out,
            y(1 to 14 - 1) => dummy127
        );


    p128_in <= x(3) & x(6) & x(10) & x(24) & x(26) & x(27) & x(40) & x(42) & x(43) & x(46) & x(52) & x(54) & x(61) & x(66) & x(68) & x(71) & x(79) & x(84) & x(87) & x(91) & x(96) & x(97) & x(100) & x(112) & x(122) & x(138) & x(146) & x(161) & x(170) & x(176) & x(179) & x(193) & x(208) & x(214) & x(215) & x(220) & x(229) & x(230) & x(233) & x(248);
    y(128) <= not(p128_out);
    p128 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111101000000011101011110111010001110011",
            TABLE => "0000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101100010101110111111000000100010101100000010001010110000000000000010001010111011110101000010001010110100001000101011110101000100001001101001100101101001011001101001100101100110100101101001100101100000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100111000100010000011100010001100001101001100101100000000000000000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p128_in,
            y(0) => p128_out,
            y(1 to 15 - 1) => dummy128
        );


    p129_in <= x(4) & x(6) & x(22) & x(37) & x(39) & x(45) & x(48) & x(52) & x(53) & x(59) & x(61) & x(65) & x(71) & x(73) & x(90) & x(114) & x(117) & x(128) & x(147) & x(156) & x(181) & x(185) & x(199) & x(203) & x(211) & x(215) & x(225) & x(227) & x(228) & x(232) & x(236) & x(243) & x(245) & x(247) & x(248);
    y(129) <= not(p129_out);
    p129 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11110010010010000011000010101100000",
            TABLE => "00000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100110001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100111101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011010000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100100010000011100010000000000010000011100011111011100010000011100010001100001110001100011100001100001110001111001110001100001110001100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 32,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p129_in,
            y(0) => p129_out,
            y(1 to 15 - 1) => dummy129
        );


    p130_in <= x(7) & x(21) & x(27) & x(34) & x(35) & x(37) & x(47) & x(50) & x(55) & x(57) & x(58) & x(61) & x(80) & x(84) & x(94) & x(98) & x(109) & x(110) & x(121) & x(122) & x(127) & x(167) & x(172) & x(177) & x(179) & x(183) & x(184) & x(189) & x(191) & x(192) & x(218) & x(222) & x(240) & x(242) & x(244) & x(248) & x(250) & x(255);
    y(130) <= not(p130_out);
    p130 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10111110100100000011001111010111110101",
            TABLE => "000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p130_in,
            y(0) => p130_out,
            y(1 to 15 - 1) => dummy130
        );


    p131_in <= x(4) & x(25) & x(31) & x(37) & x(40) & x(43) & x(45) & x(46) & x(48) & x(52) & x(72) & x(73) & x(86) & x(88) & x(95) & x(120) & x(136) & x(138) & x(157) & x(168) & x(169) & x(172) & x(177) & x(190) & x(193) & x(199) & x(218) & x(225) & x(236) & x(240) & x(250) & x(251) & x(254);
    y(131) <= not(p131_out);
    p131 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001001110101110000111100110010100",
            TABLE => "110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110100011101001011011111111",
            SHIFT => 4,
            B => 23,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p131_in,
            y(0) => p131_out,
            y(1 to 15 - 1) => dummy131
        );


    p132_in <= x(4) & x(7) & x(13) & x(18) & x(35) & x(44) & x(62) & x(68) & x(70) & x(82) & x(83) & x(85) & x(87) & x(93) & x(99) & x(107) & x(109) & x(111) & x(114) & x(132) & x(139) & x(140) & x(155) & x(168) & x(172) & x(199) & x(211) & x(221) & x(225) & x(226) & x(232) & x(235) & x(244) & x(249);
    y(132) <= not(p132_out);
    p132 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100001001000001101000111101100011",
            TABLE => "1110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101101000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010011011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010010111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101100000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010010111000100010000011100010001100001101001100101100000000000000000",
            SHIFT => 4,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p132_in,
            y(0) => p132_out,
            y(1 to 15 - 1) => dummy132
        );


    p133_in <= x(10) & x(11) & x(15) & x(27) & x(30) & x(45) & x(57) & x(59) & x(62) & x(73) & x(82) & x(83) & x(84) & x(85) & x(90) & x(92) & x(109) & x(110) & x(118) & x(128) & x(146) & x(152) & x(168) & x(169) & x(174) & x(180) & x(182) & x(189) & x(194) & x(195) & x(196) & x(200) & x(211) & x(216) & x(218) & x(225) & x(226) & x(232) & x(245) & x(253);
    y(133) <= not(p133_out);
    p133 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1011001011101011110011110000010101110011",
            TABLE => "0000100010001110000000000000100010001110111011110000100010001110000110001000111001110001000110001000111011100111000110001000111001101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010010111000100010000011100010001100001101001100101100000000000000000",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p133_in,
            y(0) => p133_out,
            y(1 to 14 - 1) => dummy133
        );


    p134_in <= x(4) & x(10) & x(14) & x(29) & x(35) & x(36) & x(57) & x(58) & x(61) & x(83) & x(87) & x(93) & x(107) & x(111) & x(114) & x(132) & x(137) & x(139) & x(140) & x(141) & x(145) & x(147) & x(156) & x(168) & x(174) & x(175) & x(179) & x(184) & x(198) & x(210) & x(213) & x(221) & x(226) & x(228) & x(235) & x(237) & x(243);
    y(134) <= not(p134_out);
    p134 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010100011110101011110001000011011101",
            TABLE => "0010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101101101010001000000010000000000000011111101110101001101010001000000110101000100001001000010001010111011110111010100110101000100001010010110011010010110100110010110011010011001011010010110011010010000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p134_in,
            y(0) => p134_out,
            y(1 to 15 - 1) => dummy134
        );


    p135_in <= x(7) & x(26) & x(30) & x(38) & x(50) & x(81) & x(87) & x(89) & x(100) & x(119) & x(132) & x(137) & x(139) & x(149) & x(156) & x(163) & x(165) & x(173) & x(174) & x(196) & x(201) & x(204) & x(212) & x(223) & x(224) & x(246) & x(252);
    y(135) <= not(p135_out);
    p135 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010110111110101100101010010",
            TABLE => "001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => 4,
            B => -32,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p135_in,
            y(0) => p135_out,
            y(1 to 14 - 1) => dummy135
        );


    p136_in <= x(6) & x(7) & x(18) & x(33) & x(35) & x(52) & x(55) & x(61) & x(62) & x(72) & x(86) & x(114) & x(118) & x(124) & x(128) & x(129) & x(137) & x(152) & x(153) & x(162) & x(165) & x(169) & x(170) & x(174) & x(181) & x(200) & x(214) & x(215) & x(223) & x(249) & x(255);
    y(136) <= not(p136_out);
    p136 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100000001001001111010100000110",
            TABLE => "1000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101101111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => 36,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p136_in,
            y(0) => p136_out,
            y(1 to 15 - 1) => dummy136
        );


    p137_in <= x(19) & x(21) & x(24) & x(29) & x(30) & x(36) & x(53) & x(56) & x(61) & x(62) & x(72) & x(80) & x(97) & x(148) & x(161) & x(175) & x(189) & x(199) & x(208) & x(216) & x(220) & x(231) & x(234) & x(248) & x(249);
    y(137) <= not(p137_out);
    p137 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000011101110000010100100",
            TABLE => "1101010001000000010000000000000011111101110101001101010001000000110101000100001001000010001010111011110111010100110101000100001010010110011010010110100110010110011010011001011010010110011010010000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101101111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101101011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p137_in,
            y(0) => p137_out,
            y(1 to 14 - 1) => dummy137
        );


    p138_in <= x(1) & x(16) & x(27) & x(30) & x(48) & x(52) & x(95) & x(99) & x(102) & x(171) & x(174) & x(175) & x(186) & x(197) & x(209) & x(221) & x(225) & x(232) & x(246) & x(250);
    y(138) <= not(p138_out);
    p138 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01000100011000000101",
            TABLE => "110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => -19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p138_in,
            y(0) => p138_out,
            y(1 to 14 - 1) => dummy138
        );


    p139_in <= x(28) & x(45) & x(54) & x(73) & x(88) & x(89) & x(120) & x(125) & x(139) & x(151) & x(158) & x(170) & x(184) & x(189) & x(198) & x(200) & x(218) & x(221) & x(225) & x(227) & x(232) & x(235) & x(240) & x(244) & x(245) & x(255);
    y(139) <= not(p139_out);
    p139 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101100101100000000111001",
            TABLE => "011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => 55,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p139_in,
            y(0) => p139_out,
            y(1 to 14 - 1) => dummy139
        );


    p140_in <= x(1) & x(7) & x(8) & x(12) & x(18) & x(21) & x(30) & x(34) & x(37) & x(42) & x(55) & x(56) & x(64) & x(65) & x(70) & x(89) & x(95) & x(101) & x(103) & x(105) & x(115) & x(127) & x(133) & x(137) & x(141) & x(151) & x(156) & x(163) & x(167) & x(177) & x(179) & x(183) & x(191) & x(194) & x(198) & x(205) & x(208) & x(214) & x(222) & x(226) & x(231) & x(240) & x(242) & x(253) & x(255);
    y(140) <= not(p140_out);
    p140 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000011100001110001010111001110001011000000010",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001101100101001011011111111",
            SHIFT => 4,
            B => 16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p140_in,
            y(0) => p140_out,
            y(1 to 15 - 1) => dummy140
        );


    p141_in <= x(4) & x(10) & x(22) & x(27) & x(31) & x(32) & x(57) & x(61) & x(66) & x(74) & x(77) & x(79) & x(111) & x(124) & x(127) & x(137) & x(142) & x(149) & x(156) & x(161) & x(162) & x(168) & x(172) & x(177) & x(184) & x(186) & x(189) & x(216) & x(228) & x(233) & x(246) & x(249) & x(253);
    y(141) <= not(p141_out);
    p141 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100000010110101001001001011010100",
            TABLE => "111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110100011101001011011111111",
            SHIFT => 4,
            B => -39,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p141_in,
            y(0) => p141_out,
            y(1 to 15 - 1) => dummy141
        );


    p142_in <= x(13) & x(19) & x(47) & x(60) & x(75) & x(87) & x(89) & x(91) & x(93) & x(99) & x(114) & x(119) & x(129) & x(135) & x(138) & x(140) & x(145) & x(151) & x(171) & x(173) & x(181) & x(186) & x(188) & x(189) & x(193) & x(197) & x(211) & x(213) & x(217) & x(226) & x(248) & x(255);
    y(142) <= not(p142_out);
    p142 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10001100110010011111100100111100",
            TABLE => "011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => 14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p142_in,
            y(0) => p142_out,
            y(1 to 15 - 1) => dummy142
        );


    p143_in <= x(8) & x(14) & x(36) & x(53) & x(61) & x(65) & x(68) & x(70) & x(87) & x(91) & x(96) & x(107) & x(115) & x(127) & x(134) & x(149) & x(155) & x(156) & x(161) & x(162) & x(165) & x(174) & x(198) & x(201) & x(203) & x(212) & x(218) & x(225) & x(226) & x(230) & x(233) & x(237) & x(240) & x(242) & x(244) & x(253);
    y(143) <= not(p143_out);
    p143 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110111111010100000110101110010111100",
            TABLE => "000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p143_in,
            y(0) => p143_out,
            y(1 to 15 - 1) => dummy143
        );


    p144_in <= x(8) & x(44) & x(46) & x(61) & x(62) & x(65) & x(66) & x(77) & x(90) & x(105) & x(116) & x(120) & x(126) & x(137) & x(140) & x(149) & x(164) & x(172) & x(198) & x(200) & x(218) & x(241) & x(246) & x(248);
    y(144) <= not(p144_out);
    p144 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101000100010111011000000",
            TABLE => "100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 5,
            B => 54,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p144_in,
            y(0) => p144_out,
            y(1 to 15 - 1) => dummy144
        );


    p145_in <= x(3) & x(16) & x(33) & x(40) & x(43) & x(54) & x(61) & x(68) & x(71) & x(78) & x(79) & x(82) & x(89) & x(119) & x(132) & x(136) & x(137) & x(149) & x(150) & x(152) & x(155) & x(156) & x(159) & x(162) & x(169) & x(173) & x(177) & x(212) & x(216) & x(231) & x(232) & x(241) & x(246);
    y(145) <= not(p145_out);
    p145 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110100011111000110011110110011000",
            TABLE => "000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 4,
            B => -29,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p145_in,
            y(0) => p145_out,
            y(1 to 15 - 1) => dummy145
        );


    p146_in <= x(3) & x(4) & x(12) & x(18) & x(27) & x(35) & x(36) & x(46) & x(61) & x(70) & x(71) & x(80) & x(85) & x(87) & x(95) & x(107) & x(109) & x(111) & x(120) & x(122) & x(124) & x(127) & x(129) & x(132) & x(135) & x(139) & x(149) & x(166) & x(168) & x(170) & x(184) & x(188) & x(191) & x(193) & x(196) & x(204) & x(206) & x(213) & x(221) & x(225) & x(226) & x(234) & x(243);
    y(146) <= not(p146_out);
    p146 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010101100110001101010001001111111011010010",
            TABLE => "1011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010010001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010011011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p146_in,
            y(0) => p146_out,
            y(1 to 15 - 1) => dummy146
        );


    p147_in <= x(7) & x(8) & x(10) & x(33) & x(35) & x(41) & x(53) & x(58) & x(79) & x(87) & x(90) & x(106) & x(115) & x(120) & x(133) & x(139) & x(141) & x(143) & x(144) & x(148) & x(156) & x(162) & x(165) & x(171) & x(172) & x(185) & x(191) & x(198) & x(201) & x(210) & x(225) & x(226) & x(230) & x(231) & x(235) & x(242) & x(244) & x(249);
    y(147) <= not(p147_out);
    p147 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10100001100101100101101010110010110011",
            TABLE => "100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 4,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p147_in,
            y(0) => p147_out,
            y(1 to 15 - 1) => dummy147
        );


    p148_in <= x(1) & x(8) & x(27) & x(31) & x(32) & x(44) & x(47) & x(55) & x(77) & x(78) & x(96) & x(99) & x(105) & x(111) & x(121) & x(127) & x(130) & x(135) & x(150) & x(177) & x(179) & x(191) & x(192) & x(195) & x(203) & x(204) & x(212) & x(214) & x(216) & x(219) & x(233) & x(238) & x(244) & x(249) & x(255);
    y(148) <= not(p148_out);
    p148 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00010100111010011100010110101011110",
            TABLE => "11011111010011010100110100000100010011010000010000000100000000001101101101001101010011010010010001001101001001000010010010110010100101100110100101101001100101100110100110010110100101100110100100101011101111110000001000101011000000100010101100000000000000100010101110111101010000100010101101000010001010111101010001000010011010011001011010010110011010011001011001101001011010011001011000010111000000010000000100000000011111110001011100010111000000010001011110000001100000011110100001111110000101110001011110000001100101100110100101101001100101100110100110010110100101100110100111011111010011010100110100000100010011010000010000000100000000001101101101001101010011010010010001001101001001000010010010110010100101100110100101101001100101100110100110010110100101100110100100100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011000000010001010110010101110111111010000100010101100101011101111011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p148_in,
            y(0) => p148_out,
            y(1 to 15 - 1) => dummy148
        );


    p149_in <= x(0) & x(10) & x(13) & x(18) & x(26) & x(28) & x(30) & x(34) & x(35) & x(36) & x(37) & x(39) & x(46) & x(52) & x(59) & x(60) & x(85) & x(102) & x(103) & x(111) & x(114) & x(129) & x(130) & x(137) & x(142) & x(151) & x(155) & x(156) & x(166) & x(174) & x(179) & x(186) & x(187) & x(196) & x(200) & x(202) & x(221) & x(243);
    y(149) <= not(p149_out);
    p149 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110110110100101101110101010010110111",
            TABLE => "000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 4,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p149_in,
            y(0) => p149_out,
            y(1 to 15 - 1) => dummy149
        );


    p150_in <= x(7) & x(38) & x(45) & x(55) & x(56) & x(75) & x(80) & x(86) & x(95) & x(102) & x(103) & x(127) & x(128) & x(139) & x(140) & x(147) & x(171) & x(189) & x(191) & x(206) & x(218) & x(220) & x(227) & x(250);
    y(150) <= not(p150_out);
    p150 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101101001010101001001110",
            TABLE => "000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 5,
            B => -26,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p150_in,
            y(0) => p150_out,
            y(1 to 15 - 1) => dummy150
        );


    p151_in <= x(8) & x(22) & x(34) & x(62) & x(68) & x(70) & x(72) & x(81) & x(87) & x(91) & x(103) & x(128) & x(129) & x(130) & x(139) & x(158) & x(164) & x(165) & x(168) & x(174) & x(186) & x(187) & x(189) & x(191) & x(193) & x(197) & x(199) & x(221) & x(223) & x(226) & x(233) & x(239);
    y(151) <= not(p151_out);
    p151 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00010001010000010110111111111001",
            TABLE => "111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => -25,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p151_in,
            y(0) => p151_out,
            y(1 to 15 - 1) => dummy151
        );


    p152_in <= x(4) & x(5) & x(11) & x(12) & x(16) & x(24) & x(45) & x(50) & x(54) & x(66) & x(77) & x(80) & x(82) & x(86) & x(88) & x(97) & x(114) & x(118) & x(120) & x(125) & x(143) & x(145) & x(157) & x(169) & x(172) & x(177) & x(184) & x(188) & x(190) & x(196) & x(200) & x(215) & x(218) & x(251) & x(255);
    y(152) <= not(p152_out);
    p152 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11010100001010010011000101011011110",
            TABLE => "00000100000000000100110100000100010011010000010011011111010011010010010010110010010011010010010001001101001001001101101101001101100101100110100101101001100101100110100110010110100101100110100111111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011010001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100101000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011000101011000000101011111100101011000000100000000000101011000000100010101101000010101111010010101101000010110101000010101101000010011010011001011010010110011010011001011001101001011010011001011000000010001010110010101110111111010000100010101100101011101111011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -30,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p152_in,
            y(0) => p152_out,
            y(1 to 15 - 1) => dummy152
        );


    p153_in <= x(10) & x(14) & x(29) & x(45) & x(53) & x(57) & x(58) & x(77) & x(84) & x(93) & x(97) & x(106) & x(120) & x(139) & x(141) & x(150) & x(158) & x(180) & x(191) & x(194) & x(195) & x(198) & x(201) & x(218) & x(225) & x(231) & x(242) & x(244) & x(245);
    y(153) <= not(p153_out);
    p153 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10100111100110010010110111011",
            TABLE => "01000000110101000000000001000000110101001111110101000000110101000100001011010100001010110100001011010100101111010100001011010100011010011001011010010110011010011001011001101001011010011001011000000000010000000100000011010100010000001101010011010100111111010010101101000010010000101101010001000010110101001101010010111101100101100110100101101001100101100110100110010110100101100110100110001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100100000100010011010000000000000100010011011101111100000100010011010010010001001101101100100010010001001101110110110010010001001101100101100110100101101001100101100110100110010110100101100110100100010000011100010111000111110111000110000111000101110001111001111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -25,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p153_in,
            y(0) => p153_out,
            y(1 to 14 - 1) => dummy153
        );


    p154_in <= x(6) & x(8) & x(53) & x(61) & x(63) & x(68) & x(72) & x(76) & x(96) & x(107) & x(108) & x(122) & x(127) & x(129) & x(139) & x(146) & x(150) & x(160) & x(168) & x(172) & x(175) & x(179) & x(189) & x(195) & x(199) & x(211) & x(234) & x(235) & x(242) & x(244) & x(246) & x(247);
    y(154) <= not(p154_out);
    p154 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00010001011110001011111010000111",
            TABLE => "111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 4,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p154_in,
            y(0) => p154_out,
            y(1 to 15 - 1) => dummy154
        );


    p155_in <= x(24) & x(38) & x(43) & x(44) & x(46) & x(50) & x(55) & x(61) & x(86) & x(98) & x(99) & x(103) & x(109) & x(117) & x(142) & x(156) & x(167) & x(170) & x(176) & x(177) & x(184) & x(193) & x(198) & x(210) & x(213) & x(214) & x(218) & x(219) & x(224) & x(237) & x(248) & x(250) & x(252);
    y(155) <= not(p155_out);
    p155 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001111001101110011001101000011011",
            TABLE => "000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001011100010110100111111111",
            SHIFT => 4,
            B => 50,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p155_in,
            y(0) => p155_out,
            y(1 to 15 - 1) => dummy155
        );


    p156_in <= x(4) & x(10) & x(14) & x(37) & x(42) & x(49) & x(53) & x(72) & x(77) & x(82) & x(83) & x(90) & x(110) & x(122) & x(128) & x(143) & x(172) & x(179) & x(196) & x(234) & x(245) & x(247) & x(255);
    y(156) <= not(p156_out);
    p156 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11000011111110000001100",
            TABLE => "10000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100100000000000000010000000100010111000000010001011100010111011111111110100010000001100000010001011110000001000101110001011101111110100101100110100101101001100101100110100110010110100101100110100111101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011010001110111011110000100010001110100011101110011100011000100011101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -44,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p156_in,
            y(0) => p156_out,
            y(1 to 14 - 1) => dummy156
        );


    p157_in <= x(2) & x(3) & x(5) & x(10) & x(25) & x(44) & x(54) & x(55) & x(60) & x(62) & x(78) & x(86) & x(91) & x(93) & x(104) & x(112) & x(114) & x(117) & x(124) & x(128) & x(138) & x(148) & x(150) & x(159) & x(165) & x(167) & x(174) & x(196) & x(203) & x(216) & x(233) & x(247);
    y(157) <= not(p157_out);
    p157 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001011111110001011011100110000",
            TABLE => "111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => -23,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p157_in,
            y(0) => p157_out,
            y(1 to 15 - 1) => dummy157
        );


    p158_in <= x(1) & x(7) & x(10) & x(11) & x(16) & x(22) & x(27) & x(36) & x(43) & x(56) & x(62) & x(65) & x(70) & x(77) & x(84) & x(98) & x(109) & x(112) & x(127) & x(130) & x(137) & x(139) & x(142) & x(145) & x(151) & x(152) & x(165) & x(168) & x(174) & x(176) & x(183) & x(204) & x(221) & x(225) & x(229) & x(232);
    y(158) <= not(p158_out);
    p158 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000111010100100001110111000011000001",
            TABLE => "011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p158_in,
            y(0) => p158_out,
            y(1 to 15 - 1) => dummy158
        );


    p159_in <= x(6) & x(7) & x(13) & x(18) & x(35) & x(48) & x(52) & x(53) & x(59) & x(62) & x(71) & x(73) & x(76) & x(79) & x(90) & x(92) & x(93) & x(109) & x(115) & x(141) & x(166) & x(168) & x(176) & x(186) & x(199) & x(211) & x(220) & x(235) & x(245);
    y(159) <= not(p159_out);
    p159 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11110100101000001000001001110",
            TABLE => "00000000000001000000010001001101000001000100110101001101110111111011001000100100001001000100110100100100010011010100110111011011011010011001011010010110011010011001011001101001011010011001011010110010111110110010000010110010001000001011001000000000001000001011001011011011001001001011001000100100101100100100110100100100100101100110100101101001100101100110100110010110100101100110100111111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011011111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011000101011101111110000001000101011001010111011110101000010001010110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p159_in,
            y(0) => p159_out,
            y(1 to 14 - 1) => dummy159
        );


    p160_in <= x(4) & x(42) & x(60) & x(61) & x(64) & x(89) & x(93) & x(95) & x(98) & x(101) & x(103) & x(121) & x(125) & x(128) & x(147) & x(168) & x(169) & x(171) & x(177) & x(183) & x(199) & x(208) & x(210) & x(225) & x(229) & x(240) & x(241) & x(248) & x(250) & x(253);
    y(160) <= not(p160_out);
    p160 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100010101100100011001011000011",
            TABLE => "101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 28,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p160_in,
            y(0) => p160_out,
            y(1 to 15 - 1) => dummy160
        );


    p161_in <= x(7) & x(11) & x(16) & x(23) & x(29) & x(31) & x(32) & x(40) & x(43) & x(49) & x(59) & x(76) & x(78) & x(79) & x(82) & x(86) & x(88) & x(89) & x(93) & x(95) & x(112) & x(116) & x(117) & x(119) & x(129) & x(134) & x(135) & x(136) & x(155) & x(162) & x(173) & x(174) & x(191) & x(199) & x(210) & x(213) & x(214) & x(218) & x(225) & x(232) & x(250);
    y(161) <= not(p161_out);
    p161 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01011100101110011110011100100101111000011",
            TABLE => "00010111000000010111111100010111000000010000000000010111000000010001011110000001011111100001011110000001111010000001011110000001100101100110100101101001100101100110100110010110100101100110100101110001111101110001000001110001000100000111000100000000000100000111000111100111000110000111000100011000011100011000111000011000011010011001011010010110011010011001011001101001011010011001011000010111000000010000000100000000011111110001011100010111000000010001011110000001100000011110100001111110000101110001011110000001100101100110100101101001100101100110100110010110100101100110100100010111000000010000000100000000011111110001011100010111000000010001011110000001100000011110100001111110000101110001011110000001100101100110100101101001100101100110100110010110100101100110100111010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100100000010001010110010101110111111000000000000001000000010001010110100001000101011001010111011110111010100010000100100001000101011100101100110100101101001100101100110100110010110100101100110100111110111011100010111000100010000111001110111000101110001000110001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p161_in,
            y(0) => p161_out,
            y(1 to 15 - 1) => dummy161
        );


    p162_in <= x(6) & x(7) & x(17) & x(20) & x(24) & x(28) & x(30) & x(36) & x(37) & x(40) & x(56) & x(61) & x(71) & x(76) & x(87) & x(89) & x(95) & x(96) & x(103) & x(104) & x(125) & x(129) & x(133) & x(137) & x(142) & x(152) & x(154) & x(156) & x(159) & x(160) & x(161) & x(165) & x(173) & x(174) & x(199) & x(201) & x(204) & x(209) & x(229) & x(231) & x(235) & x(237) & x(238) & x(244);
    y(162) <= not(p162_out);
    p162 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11100010110010101110010101000111100010111110",
            TABLE => "000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 4,
            B => 55,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p162_in,
            y(0) => p162_out,
            y(1 to 15 - 1) => dummy162
        );


    p163_in <= x(6) & x(10) & x(34) & x(38) & x(43) & x(48) & x(52) & x(53) & x(59) & x(72) & x(73) & x(79) & x(86) & x(90) & x(103) & x(106) & x(109) & x(114) & x(118) & x(141) & x(156) & x(166) & x(168) & x(169) & x(172) & x(177) & x(185) & x(190) & x(199) & x(211);
    y(163) <= not(p163_out);
    p163 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110101001100000100101000010101",
            TABLE => "000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p163_in,
            y(0) => p163_out,
            y(1 to 14 - 1) => dummy163
        );


    p164_in <= x(20) & x(21) & x(23) & x(24) & x(34) & x(38) & x(43) & x(61) & x(64) & x(71) & x(73) & x(82) & x(89) & x(93) & x(114) & x(127) & x(135) & x(142) & x(143) & x(155) & x(156) & x(167) & x(189) & x(196) & x(197) & x(202) & x(208) & x(226) & x(230) & x(231) & x(232) & x(242) & x(255);
    y(164) <= not(p164_out);
    p164 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001011110100101010101100101101111",
            TABLE => "011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 4,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p164_in,
            y(0) => p164_out,
            y(1 to 15 - 1) => dummy164
        );


    p165_in <= x(2) & x(4) & x(5) & x(6) & x(10) & x(19) & x(35) & x(45) & x(53) & x(65) & x(69) & x(70) & x(74) & x(88) & x(93) & x(102) & x(124) & x(129) & x(134) & x(138) & x(149) & x(150) & x(151) & x(157) & x(173) & x(177) & x(190) & x(203) & x(217) & x(221) & x(226) & x(236) & x(242) & x(244) & x(250);
    y(165) <= not(p165_out);
    p165 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11110000000010000010110001100000010",
            TABLE => "00000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100111101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011000001000100011100000000000001000100011101110111100001000100011100001100010001110011100010001100010001110111001110001100010001110011010011001011010010110011010011001011001101001011010011001011010000000111010001110100011111110000000001000000010000000111010001000000111101000111010000111111000010111100000011000000111101000100101100110100101101001100101100110100110010110100101100110100111111011101100101011001000100000110110111011001010110010001001000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p165_in,
            y(0) => p165_out,
            y(1 to 15 - 1) => dummy165
        );


    p166_in <= x(0) & x(2) & x(22) & x(36) & x(44) & x(65) & x(89) & x(96) & x(100) & x(103) & x(117) & x(144) & x(159) & x(162) & x(169) & x(176) & x(179) & x(189) & x(190) & x(194) & x(202) & x(204) & x(217) & x(219) & x(221) & x(227) & x(238);
    y(166) <= not(p166_out);
    p166 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111000101100101110100101000",
            TABLE => "000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 4,
            B => -24,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p166_in,
            y(0) => p166_out,
            y(1 to 14 - 1) => dummy166
        );


    p167_in <= x(6) & x(10) & x(12) & x(27) & x(29) & x(30) & x(37) & x(46) & x(52) & x(55) & x(56) & x(80) & x(87) & x(91) & x(141) & x(166) & x(170) & x(176) & x(178) & x(182) & x(193) & x(223) & x(225) & x(227) & x(233) & x(239) & x(252);
    y(167) <= not(p167_out);
    p167 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110011000000100001110011100",
            TABLE => "000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001100011101001011011111111",
            SHIFT => 4,
            B => 13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p167_in,
            y(0) => p167_out,
            y(1 to 14 - 1) => dummy167
        );


    p168_in <= x(24) & x(27) & x(34) & x(42) & x(45) & x(56) & x(70) & x(80) & x(89) & x(93) & x(96) & x(102) & x(103) & x(142) & x(148) & x(169) & x(170) & x(171) & x(179) & x(182) & x(184) & x(191) & x(202) & x(206) & x(215) & x(220) & x(229) & x(230) & x(231) & x(247);
    y(168) <= not(p168_out);
    p168 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101010110010111100011000110011",
            TABLE => "001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -37,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p168_in,
            y(0) => p168_out,
            y(1 to 15 - 1) => dummy168
        );


    p169_in <= x(1) & x(7) & x(8) & x(10) & x(29) & x(33) & x(35) & x(36) & x(46) & x(53) & x(56) & x(58) & x(70) & x(72) & x(79) & x(84) & x(95) & x(106) & x(111) & x(130) & x(140) & x(161) & x(168) & x(181) & x(184) & x(185) & x(187) & x(188) & x(192) & x(197) & x(200) & x(202) & x(211) & x(213) & x(220) & x(222) & x(225) & x(230) & x(233) & x(244) & x(249);
    y(169) <= not(p169_out);
    p169 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01011000100100111101011010010110001011111",
            TABLE => "00101011000000101011111100101011000000100000000000101011000000100010101101000010101111010010101101000010110101000010101101000010011010011001011010010110011010011001011001101001011010011001011011010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100100010111011111110000000100010111000000010001011100000000000000010001011101111110100000010001011110000001000101111110100010000001100101100110100101101001100101100110100110010110100101100110100100101011000000101011111100101011000000100000000000101011000000100010101101000010101111010010101101000010110101000010101101000010011010011001011010010110011010011001011001101001011010011001011001001101000001000000010000000000110111110100110101001101000001000100110100100100001001001011001011011011010011010100110100100100011010011001011010010110011010011001011001101001011010011001011010110010001000000010000000000000111110111011001010110010001000001011001000100100001001000100110111011011101100101011001000100100100101100110100101101001100101100110100110010110100101100110100100000001000101110001011101111111100000010001011100010111011111100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 53,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p169_in,
            y(0) => p169_out,
            y(1 to 15 - 1) => dummy169
        );


    p170_in <= x(7) & x(10) & x(11) & x(12) & x(20) & x(27) & x(34) & x(37) & x(45) & x(61) & x(65) & x(71) & x(75) & x(80) & x(105) & x(119) & x(121) & x(127) & x(138) & x(151) & x(152) & x(162) & x(169) & x(173) & x(174) & x(183) & x(192) & x(193) & x(201) & x(204) & x(212) & x(221) & x(242) & x(248) & x(252);
    y(170) <= not(p170_out);
    p170 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00100000111001110100010010001010010",
            TABLE => "11101000111111101000000011101000100000001110100000000000100000001110100001111110100000011110100010000001111010000001011110000001011010011001011010010110011010011001011001101001011010011001011000101011101111110000001000101011000000100010101100000000000000100010101110111101010000100010101101000010001010111101010001000010011010011001011010010110011010011001011001101001011010011001011000000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100111101111100011101000111000001000100011100000100000001000000000001110011110001110100011100001100010001110000110000001100001110001011010011001011010010110011010011001011001101001011010011001011010110010001000000010000000000000111110111011001010110010001000001011001000100100001001000100110111011011101100101011001000100100100101100110100101101001100101100110100110010110100101100110100110110010001000001111101110110010101100100010010011011011101100101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p170_in,
            y(0) => p170_out,
            y(1 to 15 - 1) => dummy170
        );


    p171_in <= x(27) & x(31) & x(43) & x(44) & x(46) & x(47) & x(52) & x(55) & x(58) & x(62) & x(66) & x(72) & x(86) & x(91) & x(96) & x(97) & x(98) & x(120) & x(124) & x(136) & x(143) & x(146) & x(153) & x(157) & x(168) & x(170) & x(172) & x(176) & x(179) & x(193) & x(199) & x(203) & x(206) & x(215) & x(218) & x(236) & x(238) & x(239) & x(251);
    y(171) <= not(p171_out);
    p171 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111011111110110010101001111011101001010",
            TABLE => "000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => 4,
            B => 37,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p171_in,
            y(0) => p171_out,
            y(1 to 15 - 1) => dummy171
        );


    p172_in <= x(12) & x(13) & x(25) & x(27) & x(29) & x(31) & x(32) & x(34) & x(49) & x(55) & x(58) & x(60) & x(79) & x(83) & x(87) & x(88) & x(135) & x(142) & x(153) & x(155) & x(156) & x(163) & x(170) & x(176) & x(212) & x(214) & x(215) & x(219) & x(222) & x(225) & x(227) & x(232) & x(233) & x(254);
    y(172) <= not(p172_out);
    p172 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001110000100111100001101000001110",
            TABLE => "0001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010011011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101100000001000101011010000100010101110010110011010010000000000000000",
            SHIFT => 4,
            B => 62,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p172_in,
            y(0) => p172_out,
            y(1 to 15 - 1) => dummy172
        );


    p173_in <= x(0) & x(4) & x(27) & x(29) & x(32) & x(37) & x(49) & x(52) & x(65) & x(66) & x(77) & x(90) & x(91) & x(95) & x(101) & x(105) & x(113) & x(117) & x(122) & x(141) & x(142) & x(149) & x(155) & x(163) & x(167) & x(169) & x(179) & x(181) & x(193) & x(195) & x(213) & x(227) & x(234) & x(236) & x(238) & x(241);
    y(173) <= not(p173_out);
    p173 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010100001011010101000101100101011011",
            TABLE => "100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p173_in,
            y(0) => p173_out,
            y(1 to 15 - 1) => dummy173
        );


    p174_in <= x(9) & x(22) & x(36) & x(43) & x(51) & x(61) & x(65) & x(66) & x(67) & x(77) & x(80) & x(89) & x(91) & x(93) & x(95) & x(125) & x(149) & x(156) & x(158) & x(170) & x(171) & x(174) & x(177) & x(179) & x(185) & x(189) & x(193) & x(195) & x(200) & x(203) & x(206) & x(218) & x(227) & x(232) & x(241);
    y(174) <= not(p174_out);
    p174 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001110010001111000001011011101101",
            TABLE => "11110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100110001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100100000010001010110010101110111111000000000000001000000010001010110100001000101011001010111011110111010100010000100100001000101011100101100110100101101001100101100110100110010110100101100110100111111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011000000001000000000001011100000001000101110000000101111111000101111000000111101000000101111000000100010111100000010111111000010111011010011001011010010110011010011001011001101001011010011001011001001101110111110000010001001101010011011101101100100100010011010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -50,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p174_in,
            y(0) => p174_out,
            y(1 to 15 - 1) => dummy174
        );


    p175_in <= x(10) & x(30) & x(38) & x(68) & x(69) & x(71) & x(75) & x(76) & x(79) & x(89) & x(93) & x(116) & x(133) & x(139) & x(141) & x(145) & x(156) & x(194) & x(195) & x(208) & x(211) & x(225) & x(227) & x(231);
    y(175) <= not(p175_out);
    p175 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111111001000011110111101",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p175_in,
            y(0) => p175_out,
            y(1 to 14 - 1) => dummy175
        );


    p176_in <= x(0) & x(1) & x(10) & x(17) & x(20) & x(24) & x(27) & x(35) & x(36) & x(61) & x(71) & x(72) & x(86) & x(89) & x(95) & x(106) & x(108) & x(112) & x(119) & x(121) & x(124) & x(127) & x(129) & x(134) & x(137) & x(142) & x(148) & x(154) & x(156) & x(160) & x(172) & x(187) & x(198) & x(203) & x(212) & x(235) & x(242) & x(248);
    y(176) <= not(p176_out);
    p176 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110011101110100001101110000111000110",
            TABLE => "000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 4,
            B => 49,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p176_in,
            y(0) => p176_out,
            y(1 to 15 - 1) => dummy176
        );


    p177_in <= x(4) & x(6) & x(14) & x(20) & x(40) & x(56) & x(59) & x(61) & x(63) & x(71) & x(111) & x(119) & x(120) & x(126) & x(128) & x(137) & x(139) & x(143) & x(154) & x(158) & x(160) & x(166) & x(167) & x(173) & x(174) & x(200) & x(203) & x(209) & x(212) & x(214) & x(228) & x(234) & x(235) & x(243) & x(244);
    y(177) <= not(p177_out);
    p177 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11001000110010010000110101000111100",
            TABLE => "00100000000000001011001000100000101100100010000011111011101100100010010001001101101100100010010010110010001001001101101110110010011010011001011010010110011010011001011001101001011010011001011010001110111011110000100010001110000010001000111000000000000010001000111011100111000110001000111000011000100011100111000100011000100101100110100101101001100101100110100110010110100101100110100110001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100101001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011011010100010000001111110111010100010000000000000011010100010000001101010001000010101111011101010001000010001010111101010001000010100101100110100101101001100101100110100110010110100101100110100100001000100011101000111011101111000110001000111010001110111001110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p177_in,
            y(0) => p177_out,
            y(1 to 15 - 1) => dummy177
        );


    p178_in <= x(12) & x(16) & x(24) & x(35) & x(42) & x(52) & x(72) & x(81) & x(87) & x(89) & x(93) & x(96) & x(97) & x(103) & x(108) & x(114) & x(121) & x(123) & x(128) & x(129) & x(131) & x(134) & x(142) & x(152) & x(154) & x(155) & x(156) & x(165) & x(169) & x(194) & x(202) & x(233);
    y(178) <= not(p178_out);
    p178 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00010011101100011001100100010010",
            TABLE => "111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 4,
            B => 71,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p178_in,
            y(0) => p178_out,
            y(1 to 15 - 1) => dummy178
        );


    p179_in <= x(2) & x(4) & x(10) & x(14) & x(23) & x(30) & x(33) & x(34) & x(52) & x(55) & x(61) & x(83) & x(90) & x(97) & x(102) & x(111) & x(114) & x(120) & x(138) & x(141) & x(143) & x(148) & x(152) & x(156) & x(158) & x(165) & x(172) & x(195) & x(196) & x(211) & x(213) & x(214) & x(225) & x(234) & x(236) & x(243);
    y(179) <= not(p179_out);
    p179 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111011000001001001100111010101001100",
            TABLE => "000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p179_in,
            y(0) => p179_out,
            y(1 to 15 - 1) => dummy179
        );


    p180_in <= x(6) & x(27) & x(35) & x(42) & x(70) & x(73) & x(75) & x(79) & x(104) & x(118) & x(130) & x(132) & x(138) & x(140) & x(144) & x(147) & x(192) & x(196) & x(225) & x(227) & x(236) & x(237) & x(245) & x(249);
    y(180) <= not(p180_out);
    p180 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011011101001111010111010",
            TABLE => "000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p180_in,
            y(0) => p180_out,
            y(1 to 14 - 1) => dummy180
        );


    p181_in <= x(2) & x(6) & x(21) & x(27) & x(30) & x(35) & x(44) & x(55) & x(62) & x(70) & x(75) & x(90) & x(125) & x(136) & x(144) & x(147) & x(168) & x(199) & x(225) & x(231) & x(233) & x(236) & x(242) & x(243) & x(245) & x(249);
    y(181) <= not(p181_out);
    p181 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11101010000001010001100001",
            TABLE => "000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 4,
            B => 17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p181_in,
            y(0) => p181_out,
            y(1 to 14 - 1) => dummy181
        );


    p182_in <= x(6) & x(19) & x(21) & x(27) & x(29) & x(46) & x(48) & x(55) & x(61) & x(64) & x(65) & x(66) & x(75) & x(77) & x(91) & x(96) & x(97) & x(102) & x(105) & x(114) & x(122) & x(138) & x(146) & x(156) & x(163) & x(169) & x(172) & x(179) & x(195) & x(199) & x(204) & x(212) & x(216) & x(222) & x(231) & x(241) & x(243);
    y(182) <= not(p182_out);
    p182 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010100010100101101100111000100100110",
            TABLE => "0010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101101011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010010010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101100001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010011011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010010111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -36,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p182_in,
            y(0) => p182_out,
            y(1 to 15 - 1) => dummy182
        );


    p183_in <= x(7) & x(18) & x(29) & x(38) & x(46) & x(48) & x(49) & x(53) & x(61) & x(68) & x(77) & x(81) & x(89) & x(91) & x(93) & x(105) & x(109) & x(113) & x(117) & x(119) & x(122) & x(126) & x(134) & x(135) & x(148) & x(152) & x(156) & x(162) & x(169) & x(172) & x(174) & x(178) & x(189) & x(195) & x(203) & x(209) & x(225) & x(238) & x(241) & x(245) & x(251);
    y(183) <= not(p183_out);
    p183 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01100101111010111011000100010010111101101",
            TABLE => "01000000110101001101010011111101000000000100000001000000110101000100001011010100110101001011110100101011010000100100001011010100011010011001011010010110011010011001011001101001011010011001011000000010001010110010101110111111000000000000001000000010001010110100001000101011001010111011110111010100010000100100001000101011100101100110100101101001100101100110100110010110100101100110100100000010001010110000000000000010001010111011111100000010001010110100001000101011110101000100001000101011101111010100001000101011100101100110100101101001100101100110100110010110100101100110100101000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011011101111100011101000111000001000100011100000100000001000000000001110011110001110100011100001100010001110000110000001100001110001011010011001011010010110011010011001011001101001011010011001011000000001000101110000000000000001000101110111111100000001000101111000000100010111111010001000000100010111011111101000000100010111011010011001011010010110011010011001011001101001011010011001011001001101110111110000010001001101010011011101101100100100010011010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p183_in,
            y(0) => p183_out,
            y(1 to 15 - 1) => dummy183
        );


    p184_in <= x(10) & x(27) & x(38) & x(49) & x(50) & x(58) & x(61) & x(71) & x(78) & x(87) & x(116) & x(127) & x(137) & x(143) & x(160) & x(166) & x(172) & x(175) & x(179) & x(189) & x(194) & x(195) & x(196) & x(215) & x(222) & x(231) & x(250);
    y(184) <= not(p184_out);
    p184 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111011000111001100000100001",
            TABLE => "000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110110101001001011011111111",
            SHIFT => 4,
            B => 32,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p184_in,
            y(0) => p184_out,
            y(1 to 14 - 1) => dummy184
        );


    p185_in <= x(4) & x(6) & x(16) & x(18) & x(23) & x(25) & x(29) & x(40) & x(44) & x(51) & x(61) & x(63) & x(77) & x(79) & x(80) & x(82) & x(105) & x(106) & x(115) & x(126) & x(134) & x(136) & x(148) & x(153) & x(162) & x(171) & x(174) & x(178) & x(180) & x(184) & x(187) & x(195) & x(205) & x(206) & x(208) & x(215) & x(216) & x(223) & x(225) & x(247);
    y(185) <= not(p185_out);
    p185 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010010111000111000111110001110010011101",
            TABLE => "1101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010010000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101101101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010010000010001001101001001000100110110010110011010010000000000000000",
            SHIFT => 4,
            B => -21,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p185_in,
            y(0) => p185_out,
            y(1 to 15 - 1) => dummy185
        );


    p186_in <= x(6) & x(10) & x(11) & x(21) & x(24) & x(34) & x(54) & x(66) & x(80) & x(88) & x(97) & x(101) & x(157) & x(161) & x(170) & x(174) & x(198) & x(200) & x(206) & x(210) & x(211) & x(217) & x(220) & x(227) & x(231) & x(233) & x(248) & x(249);
    y(186) <= not(p186_out);
    p186 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010001111001011001110000000",
            TABLE => "1110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010000100010001110000000000000100010001110111011110000100010001110000110001000111001110001000110001000111011100111000110001000111001101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101101110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p186_in,
            y(0) => p186_out,
            y(1 to 14 - 1) => dummy186
        );


    p187_in <= x(2) & x(6) & x(8) & x(10) & x(14) & x(34) & x(46) & x(63) & x(65) & x(68) & x(70) & x(71) & x(72) & x(73) & x(77) & x(80) & x(87) & x(90) & x(91) & x(94) & x(95) & x(96) & x(98) & x(99) & x(100) & x(102) & x(109) & x(114) & x(133) & x(138) & x(141) & x(148) & x(156) & x(166) & x(168) & x(176) & x(184) & x(186) & x(191) & x(194) & x(198) & x(199) & x(211) & x(221) & x(223) & x(226) & x(233) & x(235) & x(239);
    y(187) <= not(p187_out);
    p187 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000001010000111011100110011100111101111110110001",
            TABLE => "1111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010010010101110111111000000100010101100000010001010110000000000000010001010111011110101000010001010110100001000101011110101000100001001101001100101101001011001101001100101100110100101101001100101100000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => -40,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p187_in,
            y(0) => p187_out,
            y(1 to 15 - 1) => dummy187
        );


    p188_in <= x(3) & x(7) & x(21) & x(29) & x(37) & x(40) & x(41) & x(48) & x(50) & x(73) & x(76) & x(84) & x(86) & x(95) & x(105) & x(109) & x(114) & x(120) & x(138) & x(153) & x(157) & x(167) & x(168) & x(177) & x(181) & x(191) & x(193) & x(199) & x(205) & x(212) & x(215) & x(222) & x(228) & x(235) & x(244) & x(250);
    y(188) <= not(p188_out);
    p188 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001100101111101110001110111111000011",
            TABLE => "100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p188_in,
            y(0) => p188_out,
            y(1 to 15 - 1) => dummy188
        );


    p189_in <= x(2) & x(3) & x(14) & x(21) & x(24) & x(25) & x(33) & x(40) & x(43) & x(61) & x(86) & x(101) & x(105) & x(114) & x(115) & x(120) & x(121) & x(135) & x(136) & x(142) & x(144) & x(148) & x(149) & x(153) & x(155) & x(156) & x(158) & x(161) & x(162) & x(171) & x(174) & x(176) & x(193) & x(198) & x(199) & x(201) & x(220) & x(225) & x(231) & x(242) & x(249);
    y(189) <= not(p189_out);
    p189 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00100010111011101100101000101110101100010",
            TABLE => "11101000111111101000000011101000100000001110100000000000100000001110100001111110100000011110100010000001111010000001011110000001011010011001011010010110011010011001011001101001011010011001011000000010001010110000000000000010001010111011111100000010001010110100001000101011110101000100001000101011101111010100001000101011100101100110100101101001100101100110100110010110100101100110100100000000000100000001000001110001000100000111000101110001111101111000111000011000000110000111000100011000011100010111000111100111011010011001011010010110011010011001011001101001011010011001011010110010111110110010000010110010001000001011001000000000001000001011001011011011001001001011001000100100101100100100110100100100100101100110100101101001100101100110100110010110100101100110100101110001111101110001000001110001000100000111000100000000000100000111000111100111000110000111000100011000011100011000111000011000011010011001011010010110011010011001011001101001011010011001011000010000011100010000000000010000011100011111011100010000011100010001100001110001100011100001100001110001111001110001100001110001100101100110100101101001100101100110100110010110100101100110100111111011101100101011001000100000110110111011001010110010001001000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p189_in,
            y(0) => p189_out,
            y(1 to 15 - 1) => dummy189
        );


    p190_in <= x(5) & x(14) & x(25) & x(31) & x(39) & x(48) & x(49) & x(60) & x(71) & x(86) & x(88) & x(90) & x(92) & x(100) & x(111) & x(128) & x(132) & x(140) & x(147) & x(151) & x(164) & x(166) & x(168) & x(179) & x(194) & x(201) & x(206) & x(235) & x(247) & x(248) & x(255);
    y(190) <= not(p190_out);
    p190 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110111010000111110110011000100",
            TABLE => "0000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101101000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101101011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p190_in,
            y(0) => p190_out,
            y(1 to 15 - 1) => dummy190
        );


    p191_in <= x(4) & x(10) & x(14) & x(23) & x(27) & x(34) & x(43) & x(44) & x(53) & x(55) & x(73) & x(95) & x(114) & x(116) & x(126) & x(127) & x(128) & x(134) & x(143) & x(149) & x(157) & x(169) & x(177) & x(190) & x(193) & x(199) & x(201) & x(203) & x(216) & x(222) & x(233) & x(236) & x(247);
    y(191) <= not(p191_out);
    p191 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100100010001000101010011000001000",
            TABLE => "100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 4,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p191_in,
            y(0) => p191_out,
            y(1 to 15 - 1) => dummy191
        );


    p192_in <= x(4) & x(8) & x(14) & x(22) & x(23) & x(27) & x(28) & x(33) & x(39) & x(51) & x(54) & x(74) & x(79) & x(83) & x(92) & x(103) & x(107) & x(132) & x(139) & x(142) & x(147) & x(150) & x(156) & x(161) & x(173) & x(185) & x(187) & x(200) & x(203) & x(206) & x(211) & x(217) & x(222) & x(227) & x(235) & x(236) & x(240);
    y(192) <= not(p192_out);
    p192 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101100100110110101011100010011010100",
            TABLE => "0000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010010111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101100010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010011101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010010010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p192_in,
            y(0) => p192_out,
            y(1 to 15 - 1) => dummy192
        );


    p193_in <= x(2) & x(11) & x(17) & x(21) & x(48) & x(49) & x(53) & x(56) & x(61) & x(79) & x(82) & x(91) & x(93) & x(104) & x(105) & x(118) & x(119) & x(128) & x(134) & x(144) & x(148) & x(156) & x(162) & x(165) & x(170) & x(174) & x(175) & x(194) & x(198) & x(201) & x(203) & x(206) & x(213) & x(225) & x(235) & x(242) & x(249);
    y(193) <= not(p193_out);
    p193 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110101010001110110100100101011000110",
            TABLE => "0000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010011000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101101011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010010100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101100111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => 24,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p193_in,
            y(0) => p193_out,
            y(1 to 15 - 1) => dummy193
        );


    p194_in <= x(2) & x(5) & x(24) & x(27) & x(46) & x(47) & x(55) & x(91) & x(92) & x(100) & x(110) & x(112) & x(114) & x(118) & x(121) & x(124) & x(161) & x(169) & x(172) & x(173) & x(190) & x(196) & x(203) & x(236) & x(255);
    y(194) <= not(p194_out);
    p194 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110000011110000110010100",
            TABLE => "0000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010011111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010011011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -28,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p194_in,
            y(0) => p194_out,
            y(1 to 14 - 1) => dummy194
        );


    p195_in <= x(6) & x(24) & x(30) & x(42) & x(48) & x(53) & x(54) & x(62) & x(77) & x(114) & x(116) & x(117) & x(131) & x(154) & x(170) & x(179) & x(182) & x(185) & x(186) & x(189) & x(203) & x(205) & x(208) & x(209) & x(211) & x(212) & x(218) & x(232) & x(235) & x(236) & x(241) & x(251);
    y(195) <= not(p195_out);
    p195 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01000101111101001110110101100111",
            TABLE => "110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 4,
            B => -41,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p195_in,
            y(0) => p195_out,
            y(1 to 15 - 1) => dummy195
        );


    p196_in <= x(8) & x(18) & x(26) & x(29) & x(31) & x(37) & x(41) & x(42) & x(46) & x(49) & x(66) & x(69) & x(71) & x(73) & x(87) & x(89) & x(93) & x(99) & x(105) & x(114) & x(115) & x(134) & x(136) & x(156) & x(168) & x(194) & x(203) & x(209) & x(217) & x(222) & x(224) & x(225) & x(226) & x(227) & x(229) & x(235) & x(237) & x(247) & x(255);
    y(196) <= not(p196_out);
    p196 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101011011011101101001110010001001011101",
            TABLE => "000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110010011010110100111111111",
            SHIFT => 4,
            B => 25,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p196_in,
            y(0) => p196_out,
            y(1 to 15 - 1) => dummy196
        );


    p197_in <= x(3) & x(4) & x(8) & x(10) & x(27) & x(32) & x(34) & x(49) & x(52) & x(53) & x(72) & x(77) & x(79) & x(80) & x(83) & x(100) & x(105) & x(122) & x(127) & x(130) & x(143) & x(161) & x(168) & x(172) & x(175) & x(202) & x(210) & x(231) & x(234) & x(241) & x(247);
    y(197) <= not(p197_out);
    p197 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001111110001001010111111001001",
            TABLE => "0001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101101000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p197_in,
            y(0) => p197_out,
            y(1 to 15 - 1) => dummy197
        );


    p198_in <= x(28) & x(36) & x(46) & x(49) & x(55) & x(56) & x(61) & x(69) & x(72) & x(87) & x(96) & x(103) & x(106) & x(129) & x(145) & x(150) & x(156) & x(158) & x(173) & x(175) & x(177) & x(183) & x(185) & x(186) & x(188) & x(203) & x(209) & x(226) & x(228) & x(234) & x(247) & x(250);
    y(198) <= not(p198_out);
    p198 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00111010000110010001110111101010",
            TABLE => "001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p198_in,
            y(0) => p198_out,
            y(1 to 15 - 1) => dummy198
        );


    p199_in <= x(17) & x(23) & x(24) & x(25) & x(27) & x(29) & x(31) & x(43) & x(57) & x(86) & x(89) & x(97) & x(100) & x(105) & x(108) & x(109) & x(122) & x(123) & x(127) & x(135) & x(136) & x(137) & x(142) & x(147) & x(149) & x(153) & x(154) & x(157) & x(165) & x(167) & x(169) & x(170) & x(184) & x(187) & x(191) & x(194) & x(198) & x(203) & x(206) & x(213) & x(215) & x(220) & x(221) & x(232) & x(237) & x(243) & x(248);
    y(199) <= not(p199_out);
    p199 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10110000000110101010101011100010000011011100011",
            TABLE => "00001000100011100000000000001000100011101110111100001000100011100001100010001110011100010001100010001110111001110001100010001110011010011001011010010110011010011001011001101001011010011001011011111101110101001101010001000000110101000100000001000000000000001011110111010100110101000100001011010100010000100100001000101011011010011001011010010110011010011001011001101001011010011001011000100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011000100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011000000000100000001000000011101000100000001110100011101000111111100001011110000001100000011110100010000001111010001110100001111110011010011001011010010110011010011001011001101001011010011001011011101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011000000001000000000001011100000001000101110000000101111111000101111000000111101000000101111000000100010111100000010111111000010111011010011001011010010110011010011001011001101001011010011001011011110111011100010111000100010000111001110111000101110001000110001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p199_in,
            y(0) => p199_out,
            y(1 to 15 - 1) => dummy199
        );


    p200_in <= x(6) & x(24) & x(36) & x(37) & x(41) & x(42) & x(46) & x(53) & x(62) & x(79) & x(88) & x(105) & x(109) & x(116) & x(118) & x(128) & x(142) & x(169) & x(172) & x(176) & x(179) & x(185) & x(195) & x(197) & x(198) & x(208) & x(209) & x(218) & x(219) & x(221) & x(232) & x(235) & x(236) & x(240) & x(245) & x(252) & x(255);
    y(200) <= not(p200_out);
    p200 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001011000100011001110010100101101011",
            TABLE => "0100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101101011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010011000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010011011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010010000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 61,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p200_in,
            y(0) => p200_out,
            y(1 to 15 - 1) => dummy200
        );


    p201_in <= x(1) & x(31) & x(35) & x(66) & x(82) & x(88) & x(90) & x(91) & x(114) & x(130) & x(157) & x(165) & x(170) & x(179) & x(196) & x(200) & x(214) & x(215) & x(218) & x(225) & x(227) & x(232) & x(233) & x(237) & x(238) & x(241) & x(245) & x(251);
    y(201) <= not(p201_out);
    p201 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010101011000001111110001111",
            TABLE => "1011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010010000100010001110000000000000100010001110111011110000100010001110000110001000111001110001000110001000111011100111000110001000111001101001100101101001011001101001100101100110100101101001100101100111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 4,
            B => -20,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p201_in,
            y(0) => p201_out,
            y(1 to 14 - 1) => dummy201
        );


    p202_in <= x(6) & x(10) & x(27) & x(31) & x(35) & x(38) & x(58) & x(62) & x(69) & x(71) & x(73) & x(75) & x(90) & x(98) & x(104) & x(111) & x(125) & x(135) & x(140) & x(147) & x(152) & x(174) & x(176) & x(177) & x(187) & x(190) & x(192) & x(199) & x(201) & x(231) & x(233) & x(236) & x(244) & x(245) & x(255);
    y(202) <= not(p202_out);
    p202 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10010110110000000101011000001110101",
            TABLE => "01001101000001000000010000000000110111110100110101001101000001000100110100100100001001001011001011011011010011010100110100100100011010011001011010010110011010011001011001101001011010011001011000001000100011100000000000001000100011101110111100001000100011100001100010001110011100010001100010001110111001110001100010001110011010011001011010010110011010011001011001101001011010011001011011111101110101001101010001000000110101000100000001000000000000001011110111010100110101000100001011010100010000100100001000101011011010011001011010010110011010011001011001101001011010011001011000101011000000101011111100101011000000100000000000101011000000100010101101000010101111010010101101000010110101000010101101000010011010011001011010010110011010011001011001101001011010011001011011110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100101001101000001001101111101001101010011010010010011011011010011010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p202_in,
            y(0) => p202_out,
            y(1 to 15 - 1) => dummy202
        );


    p203_in <= x(34) & x(38) & x(51) & x(61) & x(65) & x(66) & x(67) & x(70) & x(77) & x(88) & x(119) & x(122) & x(154) & x(156) & x(157) & x(170) & x(171) & x(183) & x(185) & x(198) & x(203) & x(204) & x(209) & x(210) & x(232) & x(235) & x(248);
    y(203) <= not(p203_out);
    p203 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010001100101011111000101110",
            TABLE => "110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001001010110110100111111111",
            SHIFT => 4,
            B => 61,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p203_in,
            y(0) => p203_out,
            y(1 to 14 - 1) => dummy203
        );


    p204_in <= x(2) & x(5) & x(34) & x(46) & x(56) & x(57) & x(66) & x(97) & x(102) & x(103) & x(113) & x(116) & x(121) & x(149) & x(154) & x(161) & x(169) & x(170) & x(179) & x(189) & x(203) & x(209) & x(212) & x(215) & x(220) & x(228) & x(231) & x(232) & x(251);
    y(204) <= not(p204_out);
    p204 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00011010101011000111000001010",
            TABLE => "10111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100100100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011001000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011010000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100110110010111110110010000010110010101100101101101100100100101100101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 38,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p204_in,
            y(0) => p204_out,
            y(1 to 14 - 1) => dummy204
        );


    p205_in <= x(4) & x(5) & x(29) & x(31) & x(41) & x(42) & x(43) & x(46) & x(52) & x(59) & x(66) & x(72) & x(77) & x(82) & x(86) & x(89) & x(102) & x(128) & x(143) & x(148) & x(157) & x(170) & x(172) & x(179) & x(187) & x(193) & x(196) & x(218) & x(227) & x(232) & x(233) & x(241) & x(245) & x(246) & x(255);
    y(205) <= not(p205_out);
    p205 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00110111111000111110111101100110001",
            TABLE => "01001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011000000000000000100000001000101011000000100010101100101011101111111101010001000010010000100010101101000010001010110010101110111101011010011001011010010110011010011001011001101001011010011001011000010111011111110000000100010111000000010001011100000000000000010001011101111110100000010001011110000001000101111110100010000001100101100110100101101001100101100110100110010110100101100110100100000001000101110000000000000001000101110111111100000001000101111000000100010111111010001000000100010111011111101000000100010111011010011001011010010110011010011001011001101001011010011001011001000000110101001101010011111101000000000100000001000000110101000100001011010100110101001011110100101011010000100100001011010100011010011001011010010110011010011001011001101001011010011001011011010100010000001111110111010100110101000100001010111101110101001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 65,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p205_in,
            y(0) => p205_out,
            y(1 to 15 - 1) => dummy205
        );


    p206_in <= x(6) & x(7) & x(25) & x(33) & x(42) & x(43) & x(52) & x(53) & x(65) & x(86) & x(88) & x(93) & x(95) & x(106) & x(118) & x(120) & x(126) & x(137) & x(158) & x(165) & x(169) & x(171) & x(193) & x(198) & x(199) & x(215) & x(219) & x(220) & x(225) & x(231) & x(235) & x(242);
    y(206) <= not(p206_out);
    p206 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11100000100111110101000100111100",
            TABLE => "000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p206_in,
            y(0) => p206_out,
            y(1 to 15 - 1) => dummy206
        );


    p207_in <= x(6) & x(7) & x(11) & x(17) & x(27) & x(30) & x(36) & x(38) & x(52) & x(73) & x(76) & x(88) & x(95) & x(117) & x(156) & x(169) & x(171) & x(187) & x(197) & x(199) & x(219) & x(225) & x(238) & x(242) & x(246) & x(250) & x(254) & x(255);
    y(207) <= not(p207_out);
    p207 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010001011110101110100011100",
            TABLE => "1110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010011101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010010000100010001110000110001000111001101001100101100000000000000000",
            SHIFT => 4,
            B => -42,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p207_in,
            y(0) => p207_out,
            y(1 to 14 - 1) => dummy207
        );


    p208_in <= x(10) & x(13) & x(15) & x(48) & x(53) & x(59) & x(61) & x(73) & x(77) & x(82) & x(90) & x(92) & x(110) & x(118) & x(126) & x(141) & x(159) & x(168) & x(169) & x(187) & x(188) & x(189) & x(194) & x(196) & x(199) & x(200) & x(203) & x(211) & x(215) & x(216) & x(222) & x(244) & x(245) & x(251);
    y(208) <= not(p208_out);
    p208 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010100111111011011010001110110011",
            TABLE => "0010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010011000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100111000100010000011100010001100001101001100101100000000000000000",
            SHIFT => 4,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p208_in,
            y(0) => p208_out,
            y(1 to 15 - 1) => dummy208
        );


    p209_in <= x(18) & x(29) & x(31) & x(34) & x(42) & x(51) & x(59) & x(62) & x(75) & x(82) & x(90) & x(93) & x(102) & x(111) & x(161) & x(170) & x(177) & x(185) & x(194) & x(198) & x(208) & x(210) & x(214) & x(218) & x(232) & x(233) & x(239) & x(245);
    y(209) <= not(p209_out);
    p209 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110101000011011000011001100",
            TABLE => "0000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010011101010001000000010000000000000011111101110101001101010001000000110101000100001001000010001010111011110111010100110101000100001010010110011010010110100110010110011010011001011010010110011010010000100010001110000000000000100010001110111011110000100010001110000110001000111001110001000110001000111011100111000110001000111001101001100101101001011001101001100101100110100101101001100101101000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010000100010001110000110001000111001101001100101100000000000000000",
            SHIFT => 4,
            B => 77,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p209_in,
            y(0) => p209_out,
            y(1 to 14 - 1) => dummy209
        );


    p210_in <= x(4) & x(9) & x(22) & x(27) & x(29) & x(32) & x(43) & x(61) & x(65) & x(69) & x(70) & x(73) & x(77) & x(79) & x(93) & x(96) & x(105) & x(106) & x(112) & x(113) & x(126) & x(134) & x(136) & x(142) & x(150) & x(151) & x(156) & x(162) & x(178) & x(187) & x(190) & x(191) & x(195) & x(197) & x(208) & x(209) & x(210) & x(215) & x(225) & x(241) & x(247) & x(248);
    y(210) <= not(p210_out);
    p210 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100110111001101011000000111101111111101100",
            TABLE => "001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p210_in,
            y(0) => p210_out,
            y(1 to 15 - 1) => dummy210
        );


    p211_in <= x(7) & x(11) & x(12) & x(30) & x(34) & x(49) & x(54) & x(59) & x(65) & x(72) & x(79) & x(82) & x(83) & x(85) & x(87) & x(89) & x(93) & x(98) & x(99) & x(100) & x(124) & x(156) & x(161) & x(165) & x(174) & x(176) & x(183) & x(185) & x(189) & x(207) & x(210) & x(215) & x(217) & x(221) & x(225) & x(229) & x(254);
    y(211) <= not(p211_out);
    p211 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100001101001111100101001100011000101",
            TABLE => "1110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101100000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101100000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101000111000001000111011111000111000001000000000001000111000001000100011100001100011100111100011100001100001110001100011100001100010010110011010010110100110010110011010011001011010010110011010010100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101101011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p211_in,
            y(0) => p211_out,
            y(1 to 15 - 1) => dummy211
        );


    p212_in <= x(4) & x(8) & x(13) & x(24) & x(31) & x(34) & x(35) & x(36) & x(46) & x(56) & x(58) & x(78) & x(87) & x(93) & x(94) & x(100) & x(104) & x(107) & x(111) & x(115) & x(148) & x(156) & x(158) & x(170) & x(184) & x(185) & x(187) & x(190) & x(191) & x(193) & x(196) & x(200) & x(211) & x(213) & x(225) & x(226) & x(228) & x(235) & x(242) & x(243) & x(244) & x(248) & x(252);
    y(212) <= not(p212_out);
    p212 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000100111110010010010111100111000000000111",
            TABLE => "1111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101101101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010010111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101100001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p212_in,
            y(0) => p212_out,
            y(1 to 15 - 1) => dummy212
        );


    p213_in <= x(1) & x(4) & x(23) & x(33) & x(41) & x(56) & x(68) & x(79) & x(89) & x(137) & x(144) & x(149) & x(150) & x(152) & x(156) & x(161) & x(166) & x(172) & x(173) & x(177) & x(178) & x(180) & x(184) & x(185) & x(189) & x(203) & x(207) & x(211) & x(230) & x(231) & x(236) & x(247);
    y(213) <= not(p213_out);
    p213 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11111100101110101001000010111000",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p213_in,
            y(0) => p213_out,
            y(1 to 15 - 1) => dummy213
        );


    p214_in <= x(4) & x(8) & x(12) & x(30) & x(34) & x(42) & x(44) & x(55) & x(61) & x(70) & x(78) & x(81) & x(89) & x(98) & x(100) & x(101) & x(110) & x(127) & x(137) & x(141) & x(148) & x(156) & x(172) & x(180) & x(191) & x(198) & x(203) & x(212) & x(218) & x(223) & x(225) & x(226) & x(240) & x(244) & x(248) & x(253);
    y(214) <= not(p214_out);
    p214 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100100000011010101101110110001100101",
            TABLE => "100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p214_in,
            y(0) => p214_out,
            y(1 to 15 - 1) => dummy214
        );


    p215_in <= x(5) & x(6) & x(7) & x(10) & x(13) & x(16) & x(18) & x(22) & x(29) & x(30) & x(33) & x(34) & x(37) & x(46) & x(49) & x(53) & x(56) & x(72) & x(74) & x(79) & x(91) & x(108) & x(111) & x(120) & x(121) & x(127) & x(132) & x(148) & x(160) & x(162) & x(167) & x(173) & x(174) & x(185) & x(198) & x(204) & x(224) & x(225) & x(229) & x(231) & x(246);
    y(215) <= not(p215_out);
    p215 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000010001000011110011001100110110000001",
            TABLE => "11101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011010110010001000000010000000000000111110111011001010110010001000001011001000100100001001000100110111011011101100101011001000100100100101100110100101101001100101100110100110010110100101100110100101111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011000101011000000100000001000000000101111110010101100101011000000100010101101000010010000101101010010111101001010110010101101000010011010011001011010010110011010011001011001101001011010011001011001000000110101001101010011111101000000000100000001000000110101000100001011010100110101001011110100101011010000100100001011010100011010011001011010010110011010011001011001101001011010011001011000001000100011100000000000001000100011101110111100001000100011100001100010001110011100010001100010001110111001110001100010001110011010011001011010010110011010011001011001101001011010011001011011111101110101001101010001000000101111011101010011010100010000100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p215_in,
            y(0) => p215_out,
            y(1 to 15 - 1) => dummy215
        );


    p216_in <= x(10) & x(26) & x(27) & x(34) & x(35) & x(40) & x(41) & x(54) & x(55) & x(62) & x(64) & x(70) & x(72) & x(81) & x(83) & x(90) & x(113) & x(114) & x(124) & x(139) & x(143) & x(164) & x(165) & x(168) & x(171) & x(174) & x(192) & x(195) & x(202) & x(223) & x(225) & x(227) & x(229) & x(233) & x(236) & x(241) & x(243) & x(244) & x(245) & x(253) & x(255);
    y(216) <= not(p216_out);
    p216 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10111101110101011110101100100111101010101",
            TABLE => "00000001000101110000000000000001000101110111111100000001000101111000000100010111111010001000000100010111011111101000000100010111011010011001011010010110011010011001011001101001011010011001011000000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100100010111000000010111111100010111000000010000000000010111000000010001011110000001011111100001011110000001111010000001011110000001100101100110100101101001100101100110100110010110100101100110100100010000011100010000000000010000011100011111011100010000011100010001100001110001100011100001100001110001111001110001100001110001100101100110100101101001100101100110100110010110100101100110100111010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100100000000001000000010000010110010001000001011001010110010111110110100110100100100001001001011001000100100101100101011001011011011100101100110100101101001100101100110100110010110100101100110100101001101000001001101111101001101010011010010010011011011010011010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -37,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p216_in,
            y(0) => p216_out,
            y(1 to 15 - 1) => dummy216
        );


    p217_in <= x(4) & x(14) & x(19) & x(38) & x(44) & x(45) & x(48) & x(52) & x(59) & x(78) & x(80) & x(85) & x(88) & x(92) & x(93) & x(96) & x(101) & x(102) & x(115) & x(127) & x(133) & x(134) & x(149) & x(156) & x(161) & x(166) & x(196) & x(209) & x(225) & x(227) & x(240) & x(249);
    y(217) <= not(p217_out);
    p217 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001001000001010010010011000111",
            TABLE => "111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 4,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p217_in,
            y(0) => p217_out,
            y(1 to 15 - 1) => dummy217
        );


    p218_in <= x(0) & x(6) & x(11) & x(12) & x(15) & x(17) & x(20) & x(21) & x(30) & x(33) & x(41) & x(55) & x(72) & x(73) & x(75) & x(85) & x(92) & x(96) & x(103) & x(108) & x(114) & x(118) & x(139) & x(142) & x(155) & x(166) & x(167) & x(168) & x(169) & x(178) & x(189) & x(209) & x(215) & x(228);
    y(218) <= not(p218_out);
    p218 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110000110001001010011100010010100",
            TABLE => "1000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010011000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100010101110111111000000100010101100000010001010110000000000000010001010111011110101000010001010110100001000101011110101000100001001101001100101101001011001101001100101100110100101101001100101101101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010011000111000001000100011100001100010010110011010010000000000000000",
            SHIFT => 4,
            B => 18,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p218_in,
            y(0) => p218_out,
            y(1 to 15 - 1) => dummy218
        );


    p219_in <= x(7) & x(17) & x(19) & x(21) & x(27) & x(31) & x(53) & x(57) & x(62) & x(65) & x(91) & x(100) & x(102) & x(111) & x(114) & x(116) & x(124) & x(161) & x(175) & x(180) & x(189) & x(201) & x(204) & x(215) & x(226) & x(234) & x(239) & x(244) & x(252);
    y(219) <= not(p219_out);
    p219 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01101111010110011101010111000",
            TABLE => "00010000011100010111000111110111000000000001000000010000011100010001100001110001011100011110011110001110000110000001100001110001100101100110100101101001100101100110100110010110100101100110100100000100000000000100110100000100010011010000010011011111010011010010010010110010010011010010010001001101001001001101101101001101100101100110100101101001100101100110100110010110100101100110100100010111000000010000000100000000011111110001011100010111000000010001011110000001100000011110100001111110000101110001011110000001100101100110100101101001100101100110100110010110100101100110100101001101000001001101111101001101000001000000000001001101000001000100110100100100110110110100110100100100101100100100110100100100011010011001011010010110011010011001011001101001011010011001011010000000111010001110100011111110100000011110100011101000011111101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p219_in,
            y(0) => p219_out,
            y(1 to 14 - 1) => dummy219
        );


    p220_in <= x(10) & x(23) & x(25) & x(31) & x(33) & x(44) & x(48) & x(55) & x(57) & x(58) & x(71) & x(75) & x(78) & x(83) & x(88) & x(97) & x(102) & x(107) & x(114) & x(135) & x(140) & x(146) & x(153) & x(157) & x(170) & x(191) & x(192) & x(206) & x(212) & x(215) & x(226) & x(236) & x(241) & x(247) & x(250);
    y(220) <= not(p220_out);
    p220 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00100011001110010010101000100101010",
            TABLE => "11101000111111101000000011101000100000001110100000000000100000001110100001111110100000011110100010000001111010000001011110000001011010011001011010010110011010011001011001101001011010011001011000010000000000000111000100010000011100010001000011110111011100010001100010001110011100010001100001110001000110001110011101110001100101100110100101101001100101100110100110010110100101100110100110001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100100100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011011010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100110110010111110110010000010110010101100101101101100100100101100101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p220_in,
            y(0) => p220_out,
            y(1 to 15 - 1) => dummy220
        );


    p221_in <= x(10) & x(14) & x(31) & x(38) & x(49) & x(75) & x(76) & x(87) & x(93) & x(102) & x(103) & x(141) & x(145) & x(156) & x(176) & x(189) & x(199) & x(210) & x(211) & x(217) & x(218) & x(226) & x(227) & x(231) & x(232) & x(243) & x(246) & x(250);
    y(221) <= not(p221_out);
    p221 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100111000100001100110100110",
            TABLE => "0111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101101011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010011011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010010010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101100010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 4,
            B => -24,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p221_in,
            y(0) => p221_out,
            y(1 to 14 - 1) => dummy221
        );


    p222_in <= x(6) & x(8) & x(10) & x(35) & x(38) & x(63) & x(68) & x(69) & x(76) & x(82) & x(83) & x(87) & x(93) & x(94) & x(100) & x(102) & x(104) & x(107) & x(109) & x(129) & x(134) & x(141) & x(142) & x(152) & x(156) & x(166) & x(183) & x(184) & x(193) & x(201) & x(211) & x(218) & x(225) & x(226) & x(228) & x(229) & x(235) & x(242) & x(244) & x(248);
    y(222) <= not(p222_out);
    p222 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111111000111011100101001010011011101100",
            TABLE => "0000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010011000111000001000111011111000111000001000000000001000111000001000100011100001100011100111100011100001100001110001100011100001100010010110011010010110100110010110011010011001011010010110011010010100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010000100010001110000110001000111001101001100101100000000000000000",
            SHIFT => 4,
            B => 15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p222_in,
            y(0) => p222_out,
            y(1 to 15 - 1) => dummy222
        );


    p223_in <= x(8) & x(11) & x(18) & x(29) & x(30) & x(32) & x(55) & x(60) & x(61) & x(80) & x(83) & x(90) & x(98) & x(100) & x(109) & x(119) & x(126) & x(134) & x(147) & x(152) & x(154) & x(156) & x(169) & x(171) & x(176) & x(188) & x(189) & x(193) & x(197) & x(198) & x(199) & x(201) & x(208) & x(211) & x(216) & x(219) & x(236) & x(246) & x(252);
    y(223) <= not(p223_out);
    p223 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100001000101101011010011010100100010101",
            TABLE => "110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001010011010110100111111111",
            SHIFT => 4,
            B => 40,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p223_in,
            y(0) => p223_out,
            y(1 to 15 - 1) => dummy223
        );


    p224_in <= x(6) & x(25) & x(28) & x(46) & x(67) & x(68) & x(95) & x(96) & x(114) & x(115) & x(120) & x(142) & x(153) & x(154) & x(155) & x(156) & x(160) & x(162) & x(167) & x(172) & x(178) & x(189) & x(193) & x(197) & x(198) & x(202) & x(224) & x(225) & x(226) & x(234) & x(235) & x(238) & x(246) & x(247) & x(248) & x(255);
    y(224) <= not(p224_out);
    p224 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100111111100000111100011001111110001",
            TABLE => "000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 43,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p224_in,
            y(0) => p224_out,
            y(1 to 15 - 1) => dummy224
        );


    p225_in <= x(53) & x(55) & x(61) & x(74) & x(77) & x(83) & x(90) & x(96) & x(126) & x(149) & x(156) & x(169) & x(173) & x(177) & x(186) & x(189) & x(199) & x(208) & x(216) & x(219) & x(236) & x(241) & x(250);
    y(225) <= not(p225_out);
    p225 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01111100011001110101010",
            TABLE => "00000001000101110001011101111111000000000000000100000001000101111000000100010111000101110111111011101000100000011000000100010111011010011001011010010110011010011001011001101001011010011001011010111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100100000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100110110010111110110010000010110010101100101101101100100100101100101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p225_in,
            y(0) => p225_out,
            y(1 to 14 - 1) => dummy225
        );


    p226_in <= x(4) & x(6) & x(27) & x(48) & x(52) & x(53) & x(59) & x(69) & x(85) & x(108) & x(111) & x(115) & x(118) & x(119) & x(129) & x(131) & x(137) & x(156) & x(166) & x(168) & x(169) & x(196) & x(198) & x(200) & x(203) & x(211) & x(236) & x(241);
    y(226) <= not(p226_out);
    p226 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010110101010100001110011011",
            TABLE => "0111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101100100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101101110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101100000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010010001000001110001000110000111000110010110011010010000000000000000",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p226_in,
            y(0) => p226_out,
            y(1 to 14 - 1) => dummy226
        );


    p227_in <= x(16) & x(24) & x(27) & x(29) & x(40) & x(44) & x(62) & x(66) & x(84) & x(88) & x(106) & x(108) & x(120) & x(127) & x(145) & x(150) & x(156) & x(158) & x(163) & x(174) & x(188) & x(209) & x(225) & x(228) & x(230) & x(232) & x(241);
    y(227) <= not(p227_out);
    p227 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011100101011110110011110101",
            TABLE => "000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001010011010110100111111111",
            SHIFT => 4,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p227_in,
            y(0) => p227_out,
            y(1 to 14 - 1) => dummy227
        );


    p228_in <= x(6) & x(7) & x(13) & x(18) & x(19) & x(22) & x(23) & x(31) & x(38) & x(51) & x(56) & x(66) & x(89) & x(108) & x(113) & x(152) & x(156) & x(185) & x(189) & x(190) & x(218) & x(220) & x(227) & x(232) & x(247) & x(254);
    y(228) <= not(p228_out);
    p228 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001111101110111000000101",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p228_in,
            y(0) => p228_out,
            y(1 to 14 - 1) => dummy228
        );


    p229_in <= x(6) & x(7) & x(8) & x(11) & x(13) & x(23) & x(29) & x(30) & x(33) & x(35) & x(52) & x(55) & x(57) & x(66) & x(71) & x(89) & x(96) & x(102) & x(113) & x(157) & x(161) & x(168) & x(188) & x(192) & x(195) & x(197) & x(200) & x(207) & x(215) & x(217) & x(220) & x(226) & x(232) & x(244) & x(250);
    y(229) <= not(p229_out);
    p229 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11001011000000101000101011101110010",
            TABLE => "00100000000000001011001000100000101100100010000011111011101100100010010001001101101100100010010010110010001001001101101110110010011010011001011010010110011010011001011001101001011010011001011010000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100110110010111110110010000010110010001000001011001000000000001000001011001011011011001001001011001000100100101100100100110100100100100101100110100101101001100101100110100110010110100101100110100110110010111110110010000010110010001000001011001000000000001000001011001011011011001001001011001000100100101100100100110100100100100101100110100101101001100101100110100110010110100101100110100100000000000100000001000001110001000100000111000101110001111101111000111000011000000110000111000100011000011100010111000111100111011010011001011010010110011010011001011001101001011010011001011010110010001000001111101110110010101100100010010011011011101100101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 43,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p229_in,
            y(0) => p229_out,
            y(1 to 15 - 1) => dummy229
        );


    p230_in <= x(6) & x(17) & x(27) & x(36) & x(47) & x(52) & x(55) & x(61) & x(76) & x(83) & x(90) & x(96) & x(108) & x(110) & x(114) & x(131) & x(136) & x(160) & x(168) & x(185) & x(186) & x(189) & x(192) & x(199) & x(209) & x(211) & x(233) & x(235) & x(236) & x(239) & x(243) & x(244) & x(246) & x(247) & x(249);
    y(230) <= not(p230_out);
    p230 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11000000010101011100000001110000001",
            TABLE => "10000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100111011111010011010100110100000100010011010000010000000100000000001101101101001101010011010010010001001101001001000010010010110010100101100110100101101001100101100110100110010110100101100110100100010111000000010111111100010111000000010000000000010111000000010001011110000001011111100001011110000001111010000001011110000001100101100110100101101001100101100110100110010110100101100110100111111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100001000100011101000111011101111000000000000100000001000100011100001100010001110100011101110011101110001000110000001100010001110011010011001011010010110011010011001011001101001011010011001011011111101110101001101010001000000101111011101010011010100010000100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 48,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p230_in,
            y(0) => p230_out,
            y(1 to 15 - 1) => dummy230
        );


    p231_in <= x(0) & x(2) & x(7) & x(8) & x(29) & x(31) & x(35) & x(38) & x(49) & x(58) & x(75) & x(77) & x(82) & x(88) & x(89) & x(100) & x(102) & x(106) & x(107) & x(108) & x(119) & x(121) & x(134) & x(141) & x(147) & x(154) & x(156) & x(165) & x(168) & x(171) & x(181) & x(185) & x(191) & x(202) & x(213) & x(229) & x(234) & x(242) & x(251);
    y(231) <= not(p231_out);
    p231 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001100101010100000000111000001110111010",
            TABLE => "100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => 4,
            B => 22,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p231_in,
            y(0) => p231_out,
            y(1 to 15 - 1) => dummy231
        );


    p232_in <= x(7) & x(8) & x(16) & x(22) & x(25) & x(28) & x(31) & x(40) & x(42) & x(43) & x(46) & x(49) & x(71) & x(77) & x(83) & x(86) & x(88) & x(89) & x(105) & x(111) & x(124) & x(130) & x(135) & x(137) & x(147) & x(151) & x(153) & x(156) & x(166) & x(168) & x(174) & x(175) & x(189) & x(201) & x(210) & x(212) & x(218) & x(234) & x(235) & x(243) & x(247) & x(250) & x(255);
    y(232) <= not(p232_out);
    p232 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111001011100111111011101001111001110110011",
            TABLE => "0000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p232_in,
            y(0) => p232_out,
            y(1 to 15 - 1) => dummy232
        );


    p233_in <= x(2) & x(43) & x(50) & x(57) & x(59) & x(61) & x(70) & x(73) & x(77) & x(87) & x(107) & x(109) & x(130) & x(141) & x(142) & x(143) & x(165) & x(168) & x(170) & x(176) & x(181) & x(188) & x(199) & x(213) & x(214) & x(227) & x(234) & x(243) & x(248);
    y(233) <= not(p233_out);
    p233 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001110010001110001100110011",
            TABLE => "11110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100110001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100100001000100011101000111011101111000000000000100000001000100011100001100010001110100011101110011101110001000110000001100010001110011010011001011010010110011010011001011001101001011010011001011001000000110101001101010011111101000000000100000001000000110101000100001011010100110101001011110100101011010000100100001011010100011010011001011010010110011010011001011001101001011010011001011001110001000100001111011101110001011100010001100011100111011100010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p233_in,
            y(0) => p233_out,
            y(1 to 14 - 1) => dummy233
        );


    p234_in <= x(5) & x(8) & x(23) & x(30) & x(34) & x(38) & x(47) & x(76) & x(91) & x(95) & x(100) & x(104) & x(107) & x(119) & x(121) & x(124) & x(126) & x(127) & x(132) & x(150) & x(156) & x(160) & x(165) & x(169) & x(174) & x(178) & x(201) & x(202) & x(204) & x(215) & x(216) & x(219) & x(239) & x(252) & x(253);
    y(234) <= not(p234_out);
    p234 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10100100001101001110100111110110001",
            TABLE => "01000000110101000000000001000000110101001111110101000000110101000100001011010100001010110100001011010100101111010100001011010100011010011001011010010110011010011001011001101001011010011001011011110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100101110001000100001111011101110001000100000000000001110001000100000111000100011000111001110111000100011000100011100111000100011000011010011001011010010110011010011001011001101001011010011001011001000000110101000000000001000000110101001111110101000000110101000100001011010100001010110100001011010100101111010100001011010100011010011001011010010110011010011001011001101001011010011001011000000000000001000000010001001101000001000100110101001101110111111011001000100100001001000100110100100100010011010100110111011011011010011001011010010110011010011001011001101001011010011001011011010100010000001111110111010100110101000100001010111101110101001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p234_in,
            y(0) => p234_out,
            y(1 to 16 - 1) => dummy234
        );


    p235_in <= x(3) & x(6) & x(21) & x(48) & x(53) & x(70) & x(73) & x(88) & x(106) & x(118) & x(126) & x(127) & x(156) & x(168) & x(177) & x(192) & x(196) & x(198) & x(199) & x(211) & x(213) & x(242);
    y(235) <= not(p235_out);
    p235 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000111100100101001001",
            TABLE => "0111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101100010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101101000111000001000111011111000111000001000000000001000111000001000100011100001100011100111100011100001100001110001100011100001100010010110011010010110100110010110011010011001011010010110011010010100000011010100010000101101010001101001100101100000000000000000",
            SHIFT => 5,
            B => -22,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p235_in,
            y(0) => p235_out,
            y(1 to 15 - 1) => dummy235
        );


    p236_in <= x(6) & x(17) & x(22) & x(26) & x(58) & x(64) & x(68) & x(76) & x(81) & x(83) & x(87) & x(96) & x(98) & x(110) & x(112) & x(117) & x(125) & x(139) & x(165) & x(176) & x(184) & x(185) & x(189) & x(201) & x(223) & x(233) & x(235) & x(239) & x(244) & x(245);
    y(236) <= not(p236_out);
    p236 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000011011000100110101110100111",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -42,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p236_in,
            y(0) => p236_out,
            y(1 to 14 - 1) => dummy236
        );


    p237_in <= x(9) & x(13) & x(23) & x(34) & x(40) & x(43) & x(51) & x(53) & x(55) & x(61) & x(62) & x(65) & x(70) & x(90) & x(95) & x(99) & x(121) & x(127) & x(156) & x(163) & x(167) & x(180) & x(183) & x(185) & x(191) & x(194) & x(210) & x(214) & x(216) & x(218) & x(229) & x(230) & x(231) & x(242) & x(248) & x(253);
    y(237) <= not(p237_out);
    p237 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101001000000000001111000101010010001",
            TABLE => "010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 55,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p237_in,
            y(0) => p237_out,
            y(1 to 15 - 1) => dummy237
        );


    p238_in <= x(8) & x(12) & x(17) & x(21) & x(34) & x(37) & x(50) & x(61) & x(70) & x(71) & x(88) & x(92) & x(98) & x(117) & x(118) & x(136) & x(142) & x(156) & x(165) & x(169) & x(170) & x(172) & x(176) & x(180) & x(195) & x(210) & x(214) & x(215) & x(218) & x(232) & x(240) & x(248) & x(253) & x(255);
    y(238) <= not(p238_out);
    p238 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001001000101110011010001100010010",
            TABLE => "1110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101101011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010010000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010011000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101101011001000100000101100100010010010010110011010010000000000000000",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p238_in,
            y(0) => p238_out,
            y(1 to 15 - 1) => dummy238
        );


    p239_in <= x(6) & x(27) & x(43) & x(44) & x(46) & x(57) & x(60) & x(61) & x(70) & x(73) & x(84) & x(94) & x(95) & x(98) & x(107) & x(109) & x(114) & x(137) & x(138) & x(169) & x(177) & x(182) & x(208) & x(211) & x(212) & x(216) & x(225) & x(226) & x(236) & x(250) & x(253);
    y(239) <= not(p239_out);
    p239 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001001110001000001011110001000",
            TABLE => "1000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101101110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101100000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101101110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -30,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p239_in,
            y(0) => p239_out,
            y(1 to 15 - 1) => dummy239
        );


    p240_in <= x(5) & x(6) & x(13) & x(14) & x(17) & x(23) & x(24) & x(27) & x(34) & x(36) & x(38) & x(46) & x(52) & x(56) & x(60) & x(65) & x(66) & x(68) & x(76) & x(86) & x(91) & x(95) & x(96) & x(97) & x(98) & x(100) & x(134) & x(161) & x(170) & x(179) & x(180) & x(191) & x(197) & x(198) & x(200) & x(210) & x(215) & x(226) & x(230) & x(244) & x(248);
    y(240) <= not(p240_out);
    p240 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000101011111001011100010101101000100110",
            TABLE => "11010100010000000100000000000000111111011101010011010100010000001101010001000010010000100010101110111101110101001101010001000010100101100110100101101001100101100110100110010110100101100110100100010111000000010111111100010111000000010000000000010111000000010001011110000001011111100001011110000001111010000001011110000001100101100110100101101001100101100110100110010110100101100110100100100000000000001011001000100000101100100010000011111011101100100010010001001101101100100010010010110010001001001101101110110010011010011001011010010110011010011001011001101001011010011001011000000000100000001000000011101000100000001110100011101000111111100001011110000001100000011110100010000001111010001110100001111110011010011001011010010110011010011001011001101001011010011001011000010000011100010000000000010000011100011111011100010000011100010001100001110001100011100001100001110001111001110001100001110001100101100110100101101001100101100110100110010110100101100110100111010100010000001111110111010100010000000000000011010100010000001101010001000010101111011101010001000010001010111101010001000010100101100110100101101001100101100110100110010110100101100110100110111111001010110010101100000010101111010010101100101011010000101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p240_in,
            y(0) => p240_out,
            y(1 to 15 - 1) => dummy240
        );


    p241_in <= x(4) & x(28) & x(32) & x(37) & x(39) & x(44) & x(46) & x(51) & x(52) & x(54) & x(65) & x(66) & x(86) & x(88) & x(91) & x(117) & x(120) & x(121) & x(122) & x(125) & x(127) & x(132) & x(151) & x(156) & x(158) & x(166) & x(170) & x(172) & x(173) & x(179) & x(185) & x(189) & x(193) & x(194) & x(200) & x(202) & x(203) & x(206) & x(209) & x(218) & x(224) & x(246) & x(252) & x(255);
    y(241) <= not(p241_out);
    p241 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11001101001000011001111000001011011110110100",
            TABLE => "000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => -52,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p241_in,
            y(0) => p241_out,
            y(1 to 15 - 1) => dummy241
        );


    p242_in <= x(1) & x(34) & x(46) & x(53) & x(57) & x(69) & x(96) & x(111) & x(114) & x(116) & x(117) & x(127) & x(148) & x(150) & x(156) & x(173) & x(175) & x(177) & x(185) & x(203) & x(206) & x(212) & x(222) & x(225) & x(226) & x(227) & x(229) & x(230) & x(232) & x(236);
    y(242) <= not(p242_out);
    p242 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101000010001111011001011000110",
            TABLE => "100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p242_in,
            y(0) => p242_out,
            y(1 to 14 - 1) => dummy242
        );


    p243_in <= x(4) & x(23) & x(33) & x(34) & x(42) & x(48) & x(50) & x(55) & x(56) & x(61) & x(72) & x(85) & x(97) & x(111) & x(118) & x(142) & x(152) & x(156) & x(161) & x(165) & x(180) & x(183) & x(189) & x(195) & x(200) & x(203) & x(210) & x(214) & x(215) & x(218) & x(225) & x(226) & x(230) & x(232) & x(240) & x(242) & x(248) & x(253) & x(255);
    y(243) <= not(p243_out);
    p243 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110001101011011011010001001000101100010",
            TABLE => "010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p243_in,
            y(0) => p243_out,
            y(1 to 15 - 1) => dummy243
        );


    p244_in <= x(6) & x(8) & x(28) & x(30) & x(42) & x(55) & x(56) & x(57) & x(61) & x(62) & x(68) & x(71) & x(76) & x(77) & x(84) & x(95) & x(96) & x(125) & x(131) & x(156) & x(160) & x(161) & x(163) & x(165) & x(177) & x(186) & x(194) & x(199) & x(213) & x(220) & x(223) & x(233) & x(235) & x(236) & x(237) & x(239) & x(243) & x(244) & x(245);
    y(244) <= not(p244_out);
    p244 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110110000011000110101110000001011010000",
            TABLE => "000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 4,
            B => 75,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p244_in,
            y(0) => p244_out,
            y(1 to 15 - 1) => dummy244
        );


    p245_in <= x(3) & x(7) & x(12) & x(16) & x(18) & x(38) & x(40) & x(44) & x(49) & x(56) & x(59) & x(61) & x(79) & x(99) & x(101) & x(114) & x(119) & x(127) & x(134) & x(135) & x(156) & x(162) & x(169) & x(174) & x(180) & x(183) & x(186) & x(194) & x(200) & x(201) & x(209) & x(229) & x(231) & x(245) & x(246);
    y(245) <= not(p245_out);
    p245 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11110011100011000010001011011001110",
            TABLE => "00000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100100000000100000001000000011101000100000001110100011101000111111100001011110000001100000011110100010000001111010001110100001111110011010011001011010010110011010011001011001101001011010011001011010000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100110110010001000000010000000000000111110111011001010110010001000001011001000100100001001000100110111011011101100101011001000100100100101100110100101101001100101100110100110010110100101100110100100000010000000000010101100000010001010110000001010111111001010110100001011010100001010110100001000101011010000101011110100101011100101100110100101101001100101100110100110010110100101100110100100101011101111110000001000101011001010111011110101000010001010110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -28,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p245_in,
            y(0) => p245_out,
            y(1 to 15 - 1) => dummy245
        );


    p246_in <= x(6) & x(11) & x(12) & x(26) & x(30) & x(39) & x(46) & x(49) & x(50) & x(55) & x(56) & x(61) & x(72) & x(96) & x(102) & x(112) & x(114) & x(118) & x(141) & x(142) & x(145) & x(155) & x(156) & x(173) & x(178) & x(179) & x(183) & x(184) & x(188) & x(189) & x(192) & x(215) & x(218) & x(222) & x(226) & x(247) & x(248);
    y(246) <= not(p246_out);
    p246 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100110010101110110010111001000000100",
            TABLE => "0001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010011011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010010000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101101000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => 16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p246_in,
            y(0) => p246_out,
            y(1 to 15 - 1) => dummy246
        );


    p247_in <= x(0) & x(6) & x(7) & x(11) & x(19) & x(46) & x(53) & x(55) & x(70) & x(76) & x(93) & x(101) & x(102) & x(116) & x(118) & x(130) & x(152) & x(154) & x(161) & x(193) & x(236) & x(249) & x(252);
    y(247) <= not(p247_out);
    p247 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01100100000000111011011",
            TABLE => "01000000110101001101010011111101000000000100000001000000110101000100001011010100110101001011110100101011010000100100001011010100011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100101011101111110000001000101011000000100010101100000000000000100010101110111101010000100010101101000010001010111101010001000010011010011001011010010110011010011001011001101001011010011001011000010000011100010111000111110111000110000111000101110001111001111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 43,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p247_in,
            y(0) => p247_out,
            y(1 to 14 - 1) => dummy247
        );


    p248_in <= x(1) & x(8) & x(11) & x(16) & x(21) & x(33) & x(37) & x(40) & x(55) & x(65) & x(69) & x(91) & x(96) & x(99) & x(105) & x(114) & x(133) & x(142) & x(145) & x(152) & x(156) & x(169) & x(179) & x(195) & x(198) & x(229) & x(233) & x(238) & x(255);
    y(248) <= not(p248_out);
    p248 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11010111101101000101011001001",
            TABLE => "00000100000000000100110100000100010011010000010011011111010011010010010010110010010011010010010001001101001001001101101101001101100101100110100101101001100101100110100110010110100101100110100100000000000100000001000001110001000100000111000101110001111101111000111000011000000110000111000100011000011100010111000111100111011010011001011010010110011010011001011001101001011010011001011011010100010000001111110111010100010000000000000011010100010000001101010001000010101111011101010001000010001010111101010001000010100101100110100101101001100101100110100110010110100101100110100100101011000000101011111100101011000000100000000000101011000000100010101101000010101111010010101101000010110101000010101101000010011010011001011010010110011010011001011001101001011010011001011011010100111111010100000011010100110101001011110101000010110101001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p248_in,
            y(0) => p248_out,
            y(1 to 14 - 1) => dummy248
        );


    p249_in <= x(2) & x(6) & x(8) & x(9) & x(27) & x(41) & x(58) & x(65) & x(67) & x(68) & x(71) & x(84) & x(96) & x(98) & x(106) & x(112) & x(114) & x(130) & x(148) & x(154) & x(156) & x(173) & x(191) & x(217) & x(225) & x(236) & x(253);
    y(249) <= not(p249_out);
    p249 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000010110001011010111111111",
            TABLE => "111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 4,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p249_in,
            y(0) => p249_out,
            y(1 to 14 - 1) => dummy249
        );


    p250_in <= x(10) & x(13) & x(16) & x(19) & x(24) & x(27) & x(30) & x(34) & x(35) & x(38) & x(39) & x(40) & x(64) & x(70) & x(83) & x(90) & x(95) & x(99) & x(100) & x(101) & x(102) & x(103) & x(106) & x(109) & x(121) & x(126) & x(127) & x(129) & x(148) & x(149) & x(151) & x(156) & x(176) & x(177) & x(191) & x(192) & x(195) & x(207) & x(211) & x(218) & x(225) & x(226) & x(227) & x(236) & x(242) & x(243) & x(244) & x(245) & x(253);
    y(250) <= not(p250_out);
    p250 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110000110110101101001001001011001010101011111010",
            TABLE => "1000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101101000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101100000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -25,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p250_in,
            y(0) => p250_out,
            y(1 to 15 - 1) => dummy250
        );


    p251_in <= x(2) & x(4) & x(68) & x(73) & x(82) & x(88) & x(89) & x(90) & x(106) & x(107) & x(120) & x(125) & x(133) & x(158) & x(165) & x(167) & x(175) & x(180) & x(189) & x(200) & x(201) & x(203) & x(212) & x(218) & x(220) & x(223) & x(225) & x(230) & x(233) & x(235) & x(244) & x(245) & x(253);
    y(251) <= not(p251_out);
    p251 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101001100000010101001110000011000",
            TABLE => "010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 4,
            B => 16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p251_in,
            y(0) => p251_out,
            y(1 to 15 - 1) => dummy251
        );


    p252_in <= x(10) & x(27) & x(36) & x(44) & x(46) & x(61) & x(65) & x(66) & x(80) & x(91) & x(93) & x(94) & x(97) & x(100) & x(111) & x(121) & x(130) & x(136) & x(137) & x(145) & x(148) & x(162) & x(166) & x(170) & x(177) & x(179) & x(185) & x(189) & x(193) & x(200) & x(203) & x(204) & x(206) & x(213) & x(246) & x(252);
    y(252) <= not(p252_out);
    p252 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000101100010111010010100101101100110",
            TABLE => "110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -60,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p252_in,
            y(0) => p252_out,
            y(1 to 15 - 1) => dummy252
        );


    p253_in <= x(4) & x(6) & x(10) & x(30) & x(34) & x(53) & x(68) & x(74) & x(87) & x(90) & x(91) & x(92) & x(97) & x(108) & x(126) & x(137) & x(142) & x(143) & x(154) & x(163) & x(169) & x(172) & x(203) & x(205) & x(210) & x(211) & x(214) & x(215) & x(232) & x(235) & x(238) & x(244) & x(247) & x(248);
    y(253) <= not(p253_out);
    p253 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000110001111110111011110011000111",
            TABLE => "1111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101101000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010001011100000001000101111000000110010110011010010000000000000000",
            SHIFT => 4,
            B => -53,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p253_in,
            y(0) => p253_out,
            y(1 to 15 - 1) => dummy253
        );


    p254_in <= x(8) & x(18) & x(21) & x(27) & x(28) & x(37) & x(38) & x(42) & x(44) & x(46) & x(48) & x(52) & x(60) & x(64) & x(89) & x(92) & x(100) & x(114) & x(115) & x(117) & x(120) & x(130) & x(135) & x(141) & x(152) & x(156) & x(161) & x(165) & x(166) & x(173) & x(174) & x(178) & x(183) & x(198) & x(201) & x(206) & x(220) & x(224) & x(235) & x(242) & x(246) & x(255);
    y(254) <= not(p254_out);
    p254 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011010001010010000011000101101010100100010",
            TABLE => "001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p254_in,
            y(0) => p254_out,
            y(1 to 15 - 1) => dummy254
        );


    p255_in <= x(6) & x(10) & x(29) & x(30) & x(53) & x(56) & x(61) & x(62) & x(65) & x(72) & x(105) & x(106) & x(110) & x(114) & x(122) & x(126) & x(134) & x(135) & x(152) & x(169) & x(189) & x(195) & x(196) & x(216) & x(220) & x(221) & x(224) & x(234) & x(241) & x(248);
    y(255) <= not(p255_out);
    p255 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111100101011010001001110110011",
            TABLE => "000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p255_in,
            y(0) => p255_out,
            y(1 to 15 - 1) => dummy255
        );



end layer_2;

architecture layer_3 of layer is

    Component perceptron
    Generic (
        WEIGHTS : STD_LOGIC_VECTOR;
        SHIFT : Integer;     -- number of shift (left + or right -)
        B : Integer;          -- bias of batch norm
        BATCH_POSITIVE : Boolean    
    );
    Port ( 
        x : in STD_LOGIC_VECTOR;
        y : out STD_LOGIC_VECTOR
   );
    end component;

    -- Signals
    signal p0_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p0_out : STD_LOGIC;
	signal p1_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p1_out : STD_LOGIC;
	signal p2_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p2_out : STD_LOGIC;
	signal p3_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p3_out : STD_LOGIC;
	signal p4_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p4_out : STD_LOGIC;
	signal p5_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p5_out : STD_LOGIC;
	signal p6_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p6_out : STD_LOGIC;
	signal p7_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p7_out : STD_LOGIC;
	signal p8_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p8_out : STD_LOGIC;
	signal p9_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p9_out : STD_LOGIC;
	signal p10_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p10_out : STD_LOGIC;
	signal p11_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p11_out : STD_LOGIC;
	signal p12_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p12_out : STD_LOGIC;
	signal p13_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p13_out : STD_LOGIC;
	signal p14_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p14_out : STD_LOGIC;
	signal p15_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p15_out : STD_LOGIC;
	signal p16_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p16_out : STD_LOGIC;
	signal p17_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p17_out : STD_LOGIC;
	signal p18_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p18_out : STD_LOGIC;
	signal p19_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p19_out : STD_LOGIC;
	signal p20_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p20_out : STD_LOGIC;
	signal p21_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p21_out : STD_LOGIC;
	signal p22_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p22_out : STD_LOGIC;
	signal p23_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p23_out : STD_LOGIC;
	signal p24_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p24_out : STD_LOGIC;
	signal p25_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p25_out : STD_LOGIC;
	signal p26_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p26_out : STD_LOGIC;
	signal p27_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p27_out : STD_LOGIC;
	signal p28_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p28_out : STD_LOGIC;
	signal p29_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p29_out : STD_LOGIC;
	signal p30_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p30_out : STD_LOGIC;
	signal p31_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p31_out : STD_LOGIC;
	signal p32_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p32_out : STD_LOGIC;
	signal p33_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p33_out : STD_LOGIC;
	signal p34_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p34_out : STD_LOGIC;
	signal p35_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p35_out : STD_LOGIC;
	signal p36_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p36_out : STD_LOGIC;
	signal p37_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p37_out : STD_LOGIC;
	signal p38_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p38_out : STD_LOGIC;
	signal p39_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p39_out : STD_LOGIC;
	signal p40_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p40_out : STD_LOGIC;
	signal p41_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p41_out : STD_LOGIC;
	signal p42_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p42_out : STD_LOGIC;
	signal p43_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p43_out : STD_LOGIC;
	signal p44_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p44_out : STD_LOGIC;
	signal p45_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p45_out : STD_LOGIC;
	signal p46_in : STD_LOGIC_VECTOR(0 to 13 - 1);
	signal p46_out : STD_LOGIC;
	signal p47_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p47_out : STD_LOGIC;
	signal p48_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p48_out : STD_LOGIC;
	signal p49_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p49_out : STD_LOGIC;
	signal p50_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p50_out : STD_LOGIC;
	signal p51_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p51_out : STD_LOGIC;
	signal p52_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p52_out : STD_LOGIC;
	signal p53_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p53_out : STD_LOGIC;
	signal p54_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p54_out : STD_LOGIC;
	signal p55_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p55_out : STD_LOGIC;
	signal p56_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p56_out : STD_LOGIC;
	signal p57_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p57_out : STD_LOGIC;
	signal p58_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p58_out : STD_LOGIC;
	signal p59_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p59_out : STD_LOGIC;
	signal p60_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p60_out : STD_LOGIC;
	signal p61_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p61_out : STD_LOGIC;
	signal p62_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p62_out : STD_LOGIC;
	signal p63_in : STD_LOGIC_VECTOR(0 to 40 - 1);
	signal p63_out : STD_LOGIC;
	signal p64_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p64_out : STD_LOGIC;
	signal p65_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p65_out : STD_LOGIC;
	signal p66_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p66_out : STD_LOGIC;
	signal p67_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p67_out : STD_LOGIC;
	signal p68_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p68_out : STD_LOGIC;
	signal p69_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p69_out : STD_LOGIC;
	signal p70_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p70_out : STD_LOGIC;
	signal p71_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p71_out : STD_LOGIC;
	signal p72_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p72_out : STD_LOGIC;
	signal p73_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p73_out : STD_LOGIC;
	signal p74_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p74_out : STD_LOGIC;
	signal p75_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p75_out : STD_LOGIC;
	signal p76_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p76_out : STD_LOGIC;
	signal p77_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p77_out : STD_LOGIC;
	signal p78_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p78_out : STD_LOGIC;
	signal p79_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p79_out : STD_LOGIC;
	signal p80_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p80_out : STD_LOGIC;
	signal p81_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p81_out : STD_LOGIC;
	signal p82_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p82_out : STD_LOGIC;
	signal p83_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p83_out : STD_LOGIC;
	signal p84_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p84_out : STD_LOGIC;
	signal p85_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p85_out : STD_LOGIC;
	signal p86_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p86_out : STD_LOGIC;
	signal p87_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p87_out : STD_LOGIC;
	signal p88_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p88_out : STD_LOGIC;
	signal p89_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p89_out : STD_LOGIC;
	signal p90_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p90_out : STD_LOGIC;
	signal p91_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p91_out : STD_LOGIC;
	signal p92_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p92_out : STD_LOGIC;
	signal p93_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p93_out : STD_LOGIC;
	signal p94_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p94_out : STD_LOGIC;
	signal p95_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p95_out : STD_LOGIC;
	signal p96_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p96_out : STD_LOGIC;
	signal p97_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p97_out : STD_LOGIC;
	signal p98_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p98_out : STD_LOGIC;
	signal p99_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p99_out : STD_LOGIC;
	signal p100_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p100_out : STD_LOGIC;
	signal p101_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p101_out : STD_LOGIC;
	signal p102_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p102_out : STD_LOGIC;
	signal p103_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p103_out : STD_LOGIC;
	signal p104_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p104_out : STD_LOGIC;
	signal p105_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p105_out : STD_LOGIC;
	signal p106_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p106_out : STD_LOGIC;
	signal p107_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p107_out : STD_LOGIC;
	signal p108_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p108_out : STD_LOGIC;
	signal p109_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p109_out : STD_LOGIC;
	signal p110_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p110_out : STD_LOGIC;
	signal p111_in : STD_LOGIC_VECTOR(0 to 41 - 1);
	signal p111_out : STD_LOGIC;
	signal p112_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p112_out : STD_LOGIC;
	signal p113_in : STD_LOGIC_VECTOR(0 to 38 - 1);
	signal p113_out : STD_LOGIC;
	signal p114_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p114_out : STD_LOGIC;
	signal p115_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p115_out : STD_LOGIC;
	signal p116_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p116_out : STD_LOGIC;
	signal p117_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p117_out : STD_LOGIC;
	signal p118_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p118_out : STD_LOGIC;
	signal p119_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p119_out : STD_LOGIC;
	signal p120_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p120_out : STD_LOGIC;
	signal p121_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p121_out : STD_LOGIC;
	signal p122_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p122_out : STD_LOGIC;
	signal p123_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p123_out : STD_LOGIC;
	signal p124_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p124_out : STD_LOGIC;
	signal p125_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p125_out : STD_LOGIC;
	signal p126_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p126_out : STD_LOGIC;
	signal p127_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p127_out : STD_LOGIC;
	signal p128_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p128_out : STD_LOGIC;
	signal p129_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p129_out : STD_LOGIC;
	signal p130_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p130_out : STD_LOGIC;
	signal p131_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p131_out : STD_LOGIC;
	signal p132_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p132_out : STD_LOGIC;
	signal p133_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p133_out : STD_LOGIC;
	signal p134_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p134_out : STD_LOGIC;
	signal p135_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p135_out : STD_LOGIC;
	signal p136_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p136_out : STD_LOGIC;
	signal p137_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p137_out : STD_LOGIC;
	signal p138_in : STD_LOGIC_VECTOR(0 to 42 - 1);
	signal p138_out : STD_LOGIC;
	signal p139_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p139_out : STD_LOGIC;
	signal p140_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p140_out : STD_LOGIC;
	signal p141_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p141_out : STD_LOGIC;
	signal p142_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p142_out : STD_LOGIC;
	signal p143_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p143_out : STD_LOGIC;
	signal p144_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p144_out : STD_LOGIC;
	signal p145_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p145_out : STD_LOGIC;
	signal p146_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p146_out : STD_LOGIC;
	signal p147_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p147_out : STD_LOGIC;
	signal p148_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p148_out : STD_LOGIC;
	signal p149_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p149_out : STD_LOGIC;
	signal p150_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p150_out : STD_LOGIC;
	signal p151_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p151_out : STD_LOGIC;
	signal p152_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p152_out : STD_LOGIC;
	signal p153_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p153_out : STD_LOGIC;
	signal p154_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p154_out : STD_LOGIC;
	signal p155_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p155_out : STD_LOGIC;
	signal p156_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p156_out : STD_LOGIC;
	signal p157_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p157_out : STD_LOGIC;
	signal p158_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p158_out : STD_LOGIC;
	signal p159_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p159_out : STD_LOGIC;
	signal p160_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p160_out : STD_LOGIC;
	signal p161_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p161_out : STD_LOGIC;
	signal p162_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p162_out : STD_LOGIC;
	signal p163_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p163_out : STD_LOGIC;
	signal p164_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p164_out : STD_LOGIC;
	signal p165_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p165_out : STD_LOGIC;
	signal p166_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p166_out : STD_LOGIC;
	signal p167_in : STD_LOGIC_VECTOR(0 to 11 - 1);
	signal p167_out : STD_LOGIC;
	signal p168_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p168_out : STD_LOGIC;
	signal p169_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p169_out : STD_LOGIC;
	signal p170_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p170_out : STD_LOGIC;
	signal p171_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p171_out : STD_LOGIC;
	signal p172_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p172_out : STD_LOGIC;
	signal p173_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p173_out : STD_LOGIC;
	signal p174_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p174_out : STD_LOGIC;
	signal p175_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p175_out : STD_LOGIC;
	signal p176_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p176_out : STD_LOGIC;
	signal p177_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p177_out : STD_LOGIC;
	signal p178_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p178_out : STD_LOGIC;
	signal p179_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p179_out : STD_LOGIC;
	signal p180_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p180_out : STD_LOGIC;
	signal p181_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p181_out : STD_LOGIC;
	signal p182_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p182_out : STD_LOGIC;
	signal p183_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p183_out : STD_LOGIC;
	signal p184_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p184_out : STD_LOGIC;
	signal p185_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p185_out : STD_LOGIC;
	signal p186_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p186_out : STD_LOGIC;
	signal p187_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p187_out : STD_LOGIC;
	signal p188_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p188_out : STD_LOGIC;
	signal p189_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p189_out : STD_LOGIC;
	signal p190_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p190_out : STD_LOGIC;
	signal p191_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p191_out : STD_LOGIC;
	signal p192_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p192_out : STD_LOGIC;
	signal p193_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p193_out : STD_LOGIC;
	signal p194_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p194_out : STD_LOGIC;
	signal p195_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p195_out : STD_LOGIC;
	signal p196_in : STD_LOGIC_VECTOR(0 to 39 - 1);
	signal p196_out : STD_LOGIC;
	signal p197_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p197_out : STD_LOGIC;
	signal p198_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p198_out : STD_LOGIC;
	signal p199_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p199_out : STD_LOGIC;
	signal p200_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p200_out : STD_LOGIC;
	signal p201_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p201_out : STD_LOGIC;
	signal p202_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p202_out : STD_LOGIC;
	signal p203_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p203_out : STD_LOGIC;
	signal p204_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p204_out : STD_LOGIC;
	signal p205_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p205_out : STD_LOGIC;
	signal p206_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p206_out : STD_LOGIC;
	signal p207_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p207_out : STD_LOGIC;
	signal p208_in : STD_LOGIC_VECTOR(0 to 36 - 1);
	signal p208_out : STD_LOGIC;
	signal p209_in : STD_LOGIC_VECTOR(0 to 43 - 1);
	signal p209_out : STD_LOGIC;
	signal p210_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p210_out : STD_LOGIC;
	signal p211_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p211_out : STD_LOGIC;
	signal p212_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p212_out : STD_LOGIC;
	signal p213_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p213_out : STD_LOGIC;
	signal p214_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p214_out : STD_LOGIC;
	signal p215_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p215_out : STD_LOGIC;
	signal p216_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p216_out : STD_LOGIC;
	signal p217_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p217_out : STD_LOGIC;
	signal p218_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p218_out : STD_LOGIC;
	signal p219_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p219_out : STD_LOGIC;
	signal p220_in : STD_LOGIC_VECTOR(0 to 37 - 1);
	signal p220_out : STD_LOGIC;
	signal p221_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p221_out : STD_LOGIC;
	signal p222_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p222_out : STD_LOGIC;
	signal p223_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p223_out : STD_LOGIC;
	signal p224_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p224_out : STD_LOGIC;
	signal p225_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p225_out : STD_LOGIC;
	signal p226_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p226_out : STD_LOGIC;
	signal p227_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p227_out : STD_LOGIC;
	signal p228_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p228_out : STD_LOGIC;
	signal p229_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p229_out : STD_LOGIC;
	signal p230_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p230_out : STD_LOGIC;
	signal p231_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p231_out : STD_LOGIC;
	signal p232_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p232_out : STD_LOGIC;
	signal p233_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p233_out : STD_LOGIC;
	signal p234_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p234_out : STD_LOGIC;
	signal p235_in : STD_LOGIC_VECTOR(0 to 34 - 1);
	signal p235_out : STD_LOGIC;
	signal p236_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p236_out : STD_LOGIC;
	signal p237_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p237_out : STD_LOGIC;
	signal p238_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p238_out : STD_LOGIC;
	signal p239_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p239_out : STD_LOGIC;
	signal p240_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p240_out : STD_LOGIC;
	signal p241_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p241_out : STD_LOGIC;
	signal p242_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p242_out : STD_LOGIC;
	signal p243_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p243_out : STD_LOGIC;
	signal p244_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p244_out : STD_LOGIC;
	signal p245_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p245_out : STD_LOGIC;
	signal p246_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p246_out : STD_LOGIC;
	signal p247_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p247_out : STD_LOGIC;
	signal p248_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p248_out : STD_LOGIC;
	signal p249_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p249_out : STD_LOGIC;
	signal p250_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p250_out : STD_LOGIC;
	signal p251_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p251_out : STD_LOGIC;
	signal p252_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p252_out : STD_LOGIC;
	signal p253_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p253_out : STD_LOGIC;
	signal p254_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p254_out : STD_LOGIC;
	signal p255_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p255_out : STD_LOGIC;
	
    
    -- Dummies
    signal dummy0 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy1 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy2 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy3 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy4 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy5 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy6 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy7 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy8 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy9 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy10 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy11 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy12 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy13 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy14 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy15 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy16 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy17 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy18 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy19 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy20 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy21 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy22 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy23 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy24 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy25 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy26 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy27 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy28 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy29 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy30 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy31 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy32 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy33 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy34 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy35 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy36 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy37 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy38 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy39 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy40 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy41 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy42 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy43 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy44 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy45 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy46 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy47 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy48 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy49 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy50 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy51 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy52 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy53 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy54 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy55 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy56 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy57 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy58 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy59 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy60 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy61 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy62 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy63 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy64 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy65 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy66 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy67 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy68 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy69 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy70 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy71 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy72 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy73 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy74 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy75 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy76 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy77 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy78 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy79 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy80 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy81 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy82 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy83 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy84 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy85 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy86 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy87 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy88 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy89 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy90 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy91 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy92 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy93 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy94 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy95 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy96 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy97 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy98 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy99 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy100 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy101 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy102 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy103 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy104 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy105 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy106 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy107 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy108 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy109 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy110 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy111 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy112 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy113 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy114 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy115 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy116 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy117 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy118 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy119 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy120 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy121 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy122 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy123 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy124 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy125 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy126 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy127 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy128 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy129 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy130 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy131 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy132 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy133 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy134 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy135 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy136 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy137 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy138 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy139 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy140 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy141 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy142 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy143 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy144 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy145 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy146 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy147 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy148 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy149 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy150 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy151 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy152 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy153 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy154 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy155 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy156 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy157 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy158 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy159 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy160 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy161 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy162 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy163 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy164 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy165 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy166 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy167 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy168 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy169 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy170 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy171 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy172 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy173 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy174 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy175 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy176 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy177 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy178 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy179 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy180 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy181 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy182 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy183 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy184 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy185 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy186 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy187 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy188 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy189 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy190 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy191 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy192 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy193 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy194 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy195 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy196 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy197 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy198 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy199 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy200 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy201 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy202 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy203 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy204 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy205 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy206 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy207 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy208 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy209 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy210 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy211 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy212 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy213 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy214 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy215 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy216 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy217 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy218 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy219 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy220 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy221 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy222 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy223 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy224 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy225 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy226 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy227 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy228 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy229 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy230 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy231 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy232 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy233 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy234 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy235 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy236 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy237 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy238 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy239 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy240 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy241 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy242 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy243 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy244 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy245 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy246 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy247 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy248 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy249 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy250 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy251 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy252 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy253 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy254 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy255 : STD_LOGIC_VECTOR(0 to 13 - 2);
	 

begin

    
    p0_in <= x(7) & x(13) & x(24) & x(26) & x(38) & x(51) & x(53) & x(62) & x(69) & x(102) & x(104) & x(106) & x(109) & x(152) & x(153) & x(162) & x(166) & x(169) & x(174) & x(182) & x(185) & x(198) & x(201) & x(203) & x(207) & x(210) & x(212) & x(227) & x(229) & x(236) & x(248) & x(251) & x(252) & x(255);
    y(0) <= not(p0_out);
    p0 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010100000000000100010011010011100",
            TABLE => "1011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101101101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010010100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100000100010001110000110001000111001101001100101100000000000000000",
            SHIFT => 3,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p0_in,
            y(0) => p0_out,
            y(1 to 14 - 1) => dummy0
        );


    p1_in <= x(1) & x(4) & x(11) & x(18) & x(21) & x(29) & x(36) & x(62) & x(63) & x(77) & x(86) & x(95) & x(97) & x(100) & x(102) & x(104) & x(121) & x(122) & x(126) & x(128) & x(129) & x(131) & x(139) & x(148) & x(150) & x(156) & x(158) & x(165) & x(177) & x(179) & x(184) & x(205) & x(209) & x(229) & x(230) & x(231) & x(232) & x(233) & x(251);
    y(1) <= not(p1_out);
    p1 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010100011010100010000010100100010001011",
            TABLE => "100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001011100010110100111111111",
            SHIFT => 3,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p1_in,
            y(0) => p1_out,
            y(1 to 14 - 1) => dummy1
        );


    p2_in <= x(17) & x(28) & x(42) & x(74) & x(85) & x(89) & x(91) & x(97) & x(111) & x(116) & x(123) & x(156) & x(167) & x(177) & x(182) & x(184) & x(187) & x(190) & x(197) & x(198) & x(202) & x(214) & x(218) & x(242) & x(252);
    y(2) <= not(p2_out);
    p2 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0101101010110111100010000",
            TABLE => "0010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101100001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010010000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010011110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p2_in,
            y(0) => p2_out,
            y(1 to 14 - 1) => dummy2
        );


    p3_in <= x(14) & x(43) & x(70) & x(79) & x(95) & x(107) & x(129) & x(137) & x(140) & x(142) & x(164) & x(165) & x(179) & x(181) & x(188) & x(218) & x(232) & x(238) & x(247) & x(252);
    y(3) <= not(p3_out);
    p3 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11011000110101110111",
            TABLE => "000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 5,
            B => 19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p3_in,
            y(0) => p3_out,
            y(1 to 15 - 1) => dummy3
        );


    p4_in <= x(4) & x(6) & x(8) & x(11) & x(17) & x(27) & x(44) & x(50) & x(53) & x(62) & x(88) & x(96) & x(118) & x(119) & x(135) & x(139) & x(140) & x(143) & x(147) & x(160) & x(164) & x(172) & x(173) & x(193) & x(232) & x(251);
    y(4) <= not(p4_out);
    p4 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110010100110001011000000",
            TABLE => "000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p4_in,
            y(0) => p4_out,
            y(1 to 13 - 1) => dummy4
        );


    p5_in <= x(0) & x(16) & x(21) & x(33) & x(36) & x(45) & x(68) & x(83) & x(85) & x(103) & x(107) & x(118) & x(120) & x(121) & x(141) & x(150) & x(152) & x(174) & x(177) & x(180) & x(182) & x(186) & x(196) & x(198) & x(199) & x(202) & x(214) & x(219) & x(220) & x(232);
    y(5) <= not(p5_out);
    p5 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100101110001011111010001101010",
            TABLE => "010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p5_in,
            y(0) => p5_out,
            y(1 to 14 - 1) => dummy5
        );


    p6_in <= x(6) & x(9) & x(16) & x(48) & x(54) & x(67) & x(70) & x(72) & x(75) & x(78) & x(91) & x(95) & x(103) & x(106) & x(107) & x(113) & x(115) & x(116) & x(127) & x(137) & x(150) & x(151) & x(156) & x(164) & x(167) & x(169) & x(170) & x(172) & x(185) & x(187) & x(190) & x(196) & x(198) & x(200) & x(202) & x(210) & x(216) & x(219) & x(237) & x(252);
    y(6) <= not(p6_out);
    p6 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0101110101010101111010011101001011010011",
            TABLE => "0001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010010100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101100001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010010100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101100000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010111000100010000011100010001100001101001100101100000000000000000",
            SHIFT => 3,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p6_in,
            y(0) => p6_out,
            y(1 to 14 - 1) => dummy6
        );


    p7_in <= x(4) & x(6) & x(10) & x(18) & x(28) & x(40) & x(68) & x(85) & x(95) & x(107) & x(108) & x(112) & x(114) & x(125) & x(128) & x(152) & x(162) & x(169) & x(173) & x(205) & x(224) & x(233) & x(237) & x(244) & x(247) & x(251) & x(253);
    y(7) <= not(p7_out);
    p7 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011101110100100000010100011",
            TABLE => "000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001011100010110100111111111",
            SHIFT => 3,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p7_in,
            y(0) => p7_out,
            y(1 to 13 - 1) => dummy7
        );


    p8_in <= x(16) & x(25) & x(35) & x(41) & x(47) & x(54) & x(72) & x(73) & x(84) & x(124) & x(132) & x(133) & x(146) & x(149) & x(159) & x(165) & x(167) & x(173) & x(179) & x(190) & x(196) & x(206) & x(208) & x(217) & x(226) & x(241) & x(242) & x(254);
    y(8) <= not(p8_out);
    p8 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110100111111001000010111010",
            TABLE => "0010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101101000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101100010000010110010001001001011001001101001100101100000000000000000",
            SHIFT => 3,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p8_in,
            y(0) => p8_out,
            y(1 to 13 - 1) => dummy8
        );


    p9_in <= x(0) & x(1) & x(14) & x(16) & x(55) & x(70) & x(74) & x(86) & x(88) & x(92) & x(95) & x(103) & x(107) & x(109) & x(111) & x(112) & x(116) & x(117) & x(121) & x(130) & x(136) & x(137) & x(142) & x(156) & x(162) & x(173) & x(188) & x(190) & x(197) & x(198) & x(216) & x(219) & x(242) & x(244);
    y(9) <= not(p9_out);
    p9 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110100000100101101110101001110011",
            TABLE => "0000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101100000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010111000100010000011100010001100001101001100101100000000000000000",
            SHIFT => 3,
            B => 14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p9_in,
            y(0) => p9_out,
            y(1 to 14 - 1) => dummy9
        );


    p10_in <= x(7) & x(8) & x(25) & x(29) & x(35) & x(37) & x(53) & x(60) & x(63) & x(72) & x(75) & x(87) & x(89) & x(100) & x(133) & x(137) & x(147) & x(149) & x(153) & x(155) & x(167) & x(180) & x(186) & x(200) & x(206) & x(207) & x(215) & x(218) & x(223) & x(228) & x(233) & x(237) & x(240) & x(241) & x(254) & x(255);
    y(10) <= not(p10_out);
    p10 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110001101100100011101001100100100111",
            TABLE => "010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p10_in,
            y(0) => p10_out,
            y(1 to 14 - 1) => dummy10
        );


    p11_in <= x(4) & x(13) & x(16) & x(21) & x(52) & x(55) & x(79) & x(83) & x(99) & x(104) & x(115) & x(131) & x(135) & x(140) & x(166) & x(170) & x(172) & x(176) & x(178) & x(186) & x(189) & x(202) & x(209) & x(218) & x(220) & x(236) & x(237) & x(246) & x(248) & x(253) & x(255);
    y(11) <= not(p11_out);
    p11 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111011001110101111111110011001",
            TABLE => "0000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p11_in,
            y(0) => p11_out,
            y(1 to 15 - 1) => dummy11
        );


    p12_in <= x(12) & x(35) & x(54) & x(163) & x(179) & x(181) & x(197) & x(232) & x(246);
    y(12) <= not(p12_out);
    p12 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111110011",
            TABLE => "000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p12_in,
            y(0) => p12_out,
            y(1 to 14 - 1) => dummy12
        );


    p13_in <= x(21) & x(31) & x(41) & x(57) & x(73) & x(82) & x(89) & x(91) & x(98) & x(112) & x(132) & x(134) & x(147) & x(151) & x(154) & x(157) & x(167) & x(169) & x(184) & x(191) & x(197) & x(212) & x(221) & x(232) & x(254);
    y(13) <= not(p13_out);
    p13 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100010101010001001101010",
            TABLE => "1101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010010100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101101110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p13_in,
            y(0) => p13_out,
            y(1 to 14 - 1) => dummy13
        );


    p14_in <= x(4) & x(5) & x(10) & x(16) & x(28) & x(39) & x(40) & x(45) & x(54) & x(55) & x(62) & x(68) & x(74) & x(80) & x(99) & x(100) & x(101) & x(113) & x(124) & x(129) & x(130) & x(136) & x(140) & x(154) & x(160) & x(162) & x(175) & x(177) & x(188) & x(191) & x(195) & x(196) & x(214) & x(232) & x(234) & x(237) & x(244) & x(249) & x(250) & x(254);
    y(14) <= not(p14_out);
    p14 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0011001110011001001000111000101010110101",
            TABLE => "1000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010011000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101101011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010010001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010010100110100000100010011010010010001101001100101100000000000000000",
            SHIFT => 3,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p14_in,
            y(0) => p14_out,
            y(1 to 14 - 1) => dummy14
        );


    p15_in <= x(0) & x(1) & x(7) & x(8) & x(17) & x(18) & x(19) & x(25) & x(30) & x(39) & x(53) & x(82) & x(87) & x(91) & x(134) & x(139) & x(147) & x(153) & x(169) & x(186) & x(196) & x(206) & x(228) & x(230) & x(241) & x(251);
    y(15) <= not(p15_out);
    p15 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11110000001000001110010110",
            TABLE => "000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p15_in,
            y(0) => p15_out,
            y(1 to 13 - 1) => dummy15
        );


    p16_in <= x(0) & x(4) & x(5) & x(16) & x(33) & x(47) & x(51) & x(64) & x(84) & x(88) & x(94) & x(101) & x(107) & x(118) & x(130) & x(132) & x(149) & x(158) & x(162) & x(163) & x(170) & x(173) & x(174) & x(186) & x(188) & x(202) & x(217) & x(218) & x(219) & x(246);
    y(16) <= not(p16_out);
    p16 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111011101001011100100010001000",
            TABLE => "000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p16_in,
            y(0) => p16_out,
            y(1 to 13 - 1) => dummy16
        );


    p17_in <= x(1) & x(11) & x(29) & x(37) & x(44) & x(45) & x(46) & x(55) & x(59) & x(67) & x(75) & x(83) & x(95) & x(96) & x(108) & x(117) & x(119) & x(123) & x(126) & x(130) & x(133) & x(167) & x(168) & x(194) & x(204) & x(205) & x(208) & x(236) & x(246);
    y(17) <= not(p17_out);
    p17 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00011011000001110101000011011",
            TABLE => "10111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100110000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100100000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100111101000100000001111111011101000100000000000000011101000100000001110100010000001011111101110100010000001000101111110100010000001011010011001011010010110011010011001011001101001011010011001011000010000011100010111000111110111000110000111000101110001111001111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p17_in,
            y(0) => p17_out,
            y(1 to 13 - 1) => dummy17
        );


    p18_in <= x(3) & x(6) & x(13) & x(30) & x(34) & x(37) & x(44) & x(50) & x(55) & x(59) & x(63) & x(67) & x(69) & x(93) & x(101) & x(104) & x(121) & x(130) & x(133) & x(139) & x(144) & x(156) & x(157) & x(159) & x(188) & x(207) & x(208) & x(217) & x(221) & x(226) & x(233);
    y(18) <= not(p18_out);
    p18 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010100001011101001001001111110",
            TABLE => "1011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010011101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010010000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101101000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p18_in,
            y(0) => p18_out,
            y(1 to 14 - 1) => dummy18
        );


    p19_in <= x(4) & x(10) & x(25) & x(39) & x(53) & x(55) & x(56) & x(59) & x(77) & x(87) & x(102) & x(111) & x(122) & x(153) & x(160) & x(168) & x(169) & x(173) & x(182) & x(184) & x(207) & x(220) & x(225) & x(233) & x(240);
    y(19) <= not(p19_out);
    p19 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000100000111101111100100",
            TABLE => "1011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010011111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p19_in,
            y(0) => p19_out,
            y(1 to 14 - 1) => dummy19
        );


    p20_in <= x(6) & x(11) & x(26) & x(38) & x(49) & x(67) & x(68) & x(87) & x(95) & x(104) & x(105) & x(139) & x(144) & x(153) & x(167) & x(183) & x(195) & x(196) & x(201) & x(210) & x(238) & x(248) & x(251);
    y(20) <= not(p20_out);
    p20 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10011011000110001100011",
            TABLE => "00101011000000100000001000000000101111110010101100101011000000100010101101000010010000101101010010111101001010110010101101000010011010011001011010010110011010011001011001101001011010011001011001000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011001110001000100000001000000000000111101110111000101110001000100000111000100011000000110001000111011100111011100010111000100011000011010011001011010010110011010011001011001101001011010011001011011110111011100010111000100010000111001110111000101110001000110001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p20_in,
            y(0) => p20_out,
            y(1 to 14 - 1) => dummy20
        );


    p21_in <= x(3) & x(4) & x(6) & x(13) & x(14) & x(28) & x(30) & x(39) & x(40) & x(59) & x(62) & x(76) & x(80) & x(94) & x(124) & x(158) & x(166) & x(169) & x(173) & x(176) & x(177) & x(180) & x(192) & x(199) & x(211) & x(224) & x(238) & x(245);
    y(21) <= not(p21_out);
    p21 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010001111011111100001111000",
            TABLE => "1000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101101000000011101000100000011110100010010110011010010000000000000000",
            SHIFT => 4,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p21_in,
            y(0) => p21_out,
            y(1 to 14 - 1) => dummy21
        );


    p22_in <= x(8) & x(15) & x(19) & x(27) & x(65) & x(78) & x(79) & x(89) & x(90) & x(133) & x(134) & x(145) & x(149) & x(153) & x(166) & x(168) & x(170) & x(179) & x(189) & x(199) & x(202) & x(205) & x(209) & x(215) & x(218) & x(220) & x(230) & x(233) & x(238) & x(241) & x(245) & x(248) & x(250) & x(252) & x(255);
    y(22) <= not(p22_out);
    p22 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10001100110101110101000001100011100",
            TABLE => "01110001000100000001000000000000111101110111000101110001000100000111000100011000000110001000111011100111011100010111000100011000011010011001011010010110011010011001011001101001011010011001011001001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011000000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100111101000100000001111111011101000100000000000000011101000100000001110100010000001011111101110100010000001000101111110100010000001011010011001011010010110011010011001011001101001011010011001011010000000111010001110100011111110000000001000000010000000111010001000000111101000111010000111111000010111100000011000000111101000100101100110100101101001100101100110100110010110100101100110100100001000100011101000111011101111000110001000111010001110111001110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p22_in,
            y(0) => p22_out,
            y(1 to 15 - 1) => dummy22
        );


    p23_in <= x(1) & x(5) & x(12) & x(16) & x(20) & x(28) & x(35) & x(37) & x(47) & x(52) & x(62) & x(68) & x(72) & x(74) & x(75) & x(89) & x(113) & x(129) & x(136) & x(138) & x(143) & x(144) & x(148) & x(151) & x(156) & x(168) & x(172) & x(177) & x(182) & x(191) & x(192) & x(195) & x(204) & x(205) & x(215) & x(225) & x(232) & x(234) & x(241) & x(249) & x(251) & x(252) & x(254);
    y(23) <= not(p23_out);
    p23 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001000001111111000111100100000101100111111",
            TABLE => "1000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010011110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101100010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p23_in,
            y(0) => p23_out,
            y(1 to 14 - 1) => dummy23
        );


    p24_in <= x(4) & x(5) & x(14) & x(16) & x(22) & x(29) & x(47) & x(74) & x(76) & x(78) & x(88) & x(100) & x(107) & x(115) & x(135) & x(136) & x(148) & x(158) & x(162) & x(164) & x(170) & x(192) & x(193) & x(197) & x(202) & x(211) & x(216) & x(231) & x(232) & x(235) & x(237) & x(245);
    y(24) <= not(p24_out);
    p24 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11100010010000010010000100110101",
            TABLE => "000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 3,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p24_in,
            y(0) => p24_out,
            y(1 to 14 - 1) => dummy24
        );


    p25_in <= x(4) & x(5) & x(56) & x(72) & x(87) & x(89) & x(99) & x(107) & x(128) & x(137) & x(142) & x(161) & x(162) & x(180) & x(182) & x(206) & x(215) & x(229) & x(240) & x(245) & x(247) & x(255);
    y(25) <= not(p25_out);
    p25 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101011010101011010111",
            TABLE => "0000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101100000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010001011100000001000101111000000110010110011010010000000000000000",
            SHIFT => 4,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p25_in,
            y(0) => p25_out,
            y(1 to 14 - 1) => dummy25
        );


    p26_in <= x(9) & x(15) & x(22) & x(32) & x(33) & x(34) & x(47) & x(56) & x(63) & x(67) & x(77) & x(79) & x(91) & x(112) & x(119) & x(123) & x(128) & x(135) & x(137) & x(146) & x(149) & x(155) & x(178) & x(179) & x(183) & x(190) & x(204) & x(218) & x(232);
    y(26) <= not(p26_out);
    p26 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101101010010101111010110001",
            TABLE => "01110001111101110001000001110001000100000111000100000000000100000111000111100111000110000111000100011000011100011000111000011000011010011001011010010110011010011001011001101001011010011001011010001110000010001110111110001110000010000000000010001110000010001000111000011000111001111000111000011000011100011000111000011000100101100110100101101001100101100110100110010110100101100110100100010000011100010000000000010000011100011111011100010000011100010001100001110001100011100001100001110001111001110001100001110001100101100110100101101001100101100110100110010110100101100110100100000100000000000100110100000100010011010000010011011111010011010010010010110010010011010010010001001101001001001101101101001101100101100110100101101001100101100110100110010110100101100110100111010100010000001111110111010100110101000100001010111101110101001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p26_in,
            y(0) => p26_out,
            y(1 to 13 - 1) => dummy26
        );


    p27_in <= x(2) & x(4) & x(14) & x(15) & x(16) & x(26) & x(27) & x(34) & x(40) & x(41) & x(57) & x(64) & x(72) & x(77) & x(80) & x(101) & x(107) & x(111) & x(117) & x(130) & x(136) & x(140) & x(149) & x(161) & x(162) & x(165) & x(184) & x(187) & x(188) & x(189) & x(193) & x(196) & x(197) & x(235) & x(241) & x(244) & x(247) & x(250);
    y(27) <= not(p27_out);
    p27 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11100100000011110001100011000001110111",
            TABLE => "000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 3,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p27_in,
            y(0) => p27_out,
            y(1 to 14 - 1) => dummy27
        );


    p28_in <= x(11) & x(20) & x(46) & x(48) & x(70) & x(77) & x(79) & x(81) & x(88) & x(89) & x(92) & x(95) & x(98) & x(107) & x(109) & x(110) & x(112) & x(121) & x(131) & x(137) & x(139) & x(142) & x(145) & x(150) & x(175) & x(180) & x(188) & x(208) & x(216) & x(218) & x(229) & x(237) & x(247) & x(248) & x(251) & x(252) & x(255);
    y(28) <= not(p28_out);
    p28 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101011101010011101001101010011110011",
            TABLE => "0000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010010101110111111000000100010101100000010001010110000000000000010001010111011110101000010001010110100001000101011110101000100001001101001100101101001011001101001100101100110100101101001100101100010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 22,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p28_in,
            y(0) => p28_out,
            y(1 to 15 - 1) => dummy28
        );


    p29_in <= x(0) & x(2) & x(8) & x(9) & x(19) & x(37) & x(38) & x(43) & x(50) & x(64) & x(96) & x(101) & x(112) & x(129) & x(130) & x(131) & x(133) & x(134) & x(142) & x(188) & x(189) & x(198) & x(212) & x(218) & x(220) & x(222) & x(234) & x(246) & x(248) & x(252);
    y(29) <= not(p29_out);
    p29 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000110001100100101111001011101",
            TABLE => "101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p29_in,
            y(0) => p29_out,
            y(1 to 13 - 1) => dummy29
        );


    p30_in <= x(14) & x(26) & x(36) & x(37) & x(54) & x(57) & x(59) & x(61) & x(66) & x(86) & x(100) & x(111) & x(122) & x(147) & x(153) & x(161) & x(163) & x(165) & x(169) & x(174) & x(177) & x(179) & x(198) & x(236) & x(243) & x(254) & x(255);
    y(30) <= not(p30_out);
    p30 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001011100111011110000101110",
            TABLE => "011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001001010110110100111111111",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p30_in,
            y(0) => p30_out,
            y(1 to 14 - 1) => dummy30
        );


    p31_in <= x(0) & x(5) & x(10) & x(14) & x(16) & x(20) & x(51) & x(73) & x(74) & x(76) & x(101) & x(114) & x(118) & x(130) & x(133) & x(144) & x(152) & x(158) & x(162) & x(163) & x(166) & x(170) & x(176) & x(197) & x(211) & x(217) & x(219) & x(226) & x(239) & x(247);
    y(31) <= not(p31_out);
    p31 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110101110010111010100011010101",
            TABLE => "000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p31_in,
            y(0) => p31_out,
            y(1 to 13 - 1) => dummy31
        );


    p32_in <= x(3) & x(10) & x(29) & x(30) & x(37) & x(40) & x(45) & x(50) & x(61) & x(63) & x(66) & x(75) & x(95) & x(100) & x(131) & x(148) & x(155) & x(160) & x(164) & x(188) & x(196) & x(207) & x(209) & x(216) & x(237) & x(240);
    y(32) <= not(p32_out);
    p32 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10011001111000000010100100",
            TABLE => "001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p32_in,
            y(0) => p32_out,
            y(1 to 14 - 1) => dummy32
        );


    p33_in <= x(12) & x(26) & x(37) & x(38) & x(44) & x(50) & x(56) & x(61) & x(62) & x(71) & x(72) & x(87) & x(89) & x(103) & x(127) & x(133) & x(137) & x(142) & x(146) & x(151) & x(167) & x(170) & x(182) & x(195) & x(197) & x(205) & x(212) & x(222) & x(223) & x(248) & x(252) & x(255);
    y(33) <= not(p33_out);
    p33 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10011010000100011011000100101100",
            TABLE => "001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 4,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p33_in,
            y(0) => p33_out,
            y(1 to 15 - 1) => dummy33
        );


    p34_in <= x(19) & x(21) & x(23) & x(32) & x(35) & x(52) & x(56) & x(57) & x(59) & x(62) & x(69) & x(71) & x(76) & x(85) & x(89) & x(94) & x(113) & x(119) & x(124) & x(129) & x(142) & x(147) & x(149) & x(160) & x(172) & x(180) & x(192) & x(195) & x(197) & x(205) & x(212) & x(222) & x(229) & x(232) & x(234) & x(240) & x(241) & x(244) & x(246) & x(251) & x(252) & x(254);
    y(34) <= not(p34_out);
    p34 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000110101000100010110001111000100101010000",
            TABLE => "101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p34_in,
            y(0) => p34_out,
            y(1 to 14 - 1) => dummy34
        );


    p35_in <= x(2) & x(4) & x(13) & x(24) & x(32) & x(38) & x(44) & x(55) & x(59) & x(67) & x(69) & x(73) & x(75) & x(87) & x(104) & x(115) & x(119) & x(134) & x(141) & x(144) & x(167) & x(170) & x(171) & x(174) & x(183) & x(201) & x(203) & x(207) & x(210) & x(212) & x(222) & x(223) & x(234) & x(235) & x(240) & x(241) & x(248) & x(252);
    y(35) <= not(p35_out);
    p35 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10011111100111000001001000110101011010",
            TABLE => "000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 3,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p35_in,
            y(0) => p35_out,
            y(1 to 14 - 1) => dummy35
        );


    p36_in <= x(13) & x(17) & x(22) & x(26) & x(28) & x(33) & x(48) & x(60) & x(63) & x(64) & x(67) & x(76) & x(81) & x(84) & x(108) & x(109) & x(117) & x(124) & x(127) & x(142) & x(145) & x(149) & x(154) & x(163) & x(164) & x(165) & x(170) & x(192) & x(198) & x(216) & x(254);
    y(36) <= not(p36_out);
    p36 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111011100111101011000101111100",
            TABLE => "0000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010010000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010011011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010010000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p36_in,
            y(0) => p36_out,
            y(1 to 14 - 1) => dummy36
        );


    p37_in <= x(17) & x(25) & x(35) & x(53) & x(67) & x(68) & x(80) & x(85) & x(99) & x(101) & x(117) & x(128) & x(137) & x(156) & x(161) & x(162) & x(163) & x(172) & x(177) & x(180) & x(181) & x(186) & x(189) & x(191) & x(193) & x(194) & x(206) & x(209) & x(226) & x(230) & x(245) & x(247);
    y(37) <= not(p37_out);
    p37 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00010011110101011010100101100111",
            TABLE => "111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 3,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p37_in,
            y(0) => p37_out,
            y(1 to 14 - 1) => dummy37
        );


    p38_in <= x(4) & x(5) & x(10) & x(22) & x(32) & x(33) & x(46) & x(56) & x(73) & x(77) & x(79) & x(83) & x(91) & x(100) & x(107) & x(114) & x(119) & x(121) & x(123) & x(131) & x(135) & x(151) & x(161) & x(162) & x(166) & x(168) & x(177) & x(178) & x(194) & x(204) & x(231) & x(245);
    y(38) <= not(p38_out);
    p38 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00110101000111111100101011001000",
            TABLE => "010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 4,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p38_in,
            y(0) => p38_out,
            y(1 to 15 - 1) => dummy38
        );


    p39_in <= x(1) & x(3) & x(25) & x(44) & x(53) & x(86) & x(88) & x(99) & x(101) & x(117) & x(122) & x(129) & x(136) & x(169) & x(180) & x(188) & x(189) & x(193) & x(194) & x(203) & x(206) & x(228) & x(230) & x(236) & x(242) & x(244) & x(247) & x(254) & x(255);
    y(39) <= not(p39_out);
    p39 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00100110010000111101010110000",
            TABLE => "11010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100110001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100100010111011111110000000100010111000000010001011100000000000000010001011101111110100000010001011110000001000101111110100010000001100101100110100101101001100101100110100110010110100101100110100101001101000001001101111101001101000001000000000001001101000001000100110100100100110110110100110100100100101100100100110100100100011010011001011010010110011010011001011001101001011010011001011011101000100000001111111011101000111010001000000101111110111010000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p39_in,
            y(0) => p39_out,
            y(1 to 14 - 1) => dummy39
        );


    p40_in <= x(6) & x(8) & x(39) & x(42) & x(69) & x(70) & x(83) & x(91) & x(103) & x(105) & x(115) & x(134) & x(135) & x(151) & x(152) & x(155) & x(164) & x(171) & x(183) & x(187) & x(188) & x(193) & x(194) & x(211) & x(222) & x(234) & x(239) & x(248) & x(249) & x(252);
    y(40) <= not(p40_out);
    p40 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110001001100010101011000000110",
            TABLE => "010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p40_in,
            y(0) => p40_out,
            y(1 to 14 - 1) => dummy40
        );


    p41_in <= x(8) & x(11) & x(25) & x(26) & x(29) & x(37) & x(60) & x(63) & x(67) & x(74) & x(84) & x(90) & x(93) & x(121) & x(131) & x(140) & x(160) & x(163) & x(172) & x(175) & x(176) & x(186) & x(206) & x(209) & x(217) & x(226) & x(244);
    y(41) <= not(p41_out);
    p41 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100001010000010001000010000",
            TABLE => "110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 3,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p41_in,
            y(0) => p41_out,
            y(1 to 13 - 1) => dummy41
        );


    p42_in <= x(39) & x(44) & x(58) & x(68) & x(70) & x(86) & x(95) & x(98) & x(101) & x(103) & x(113) & x(115) & x(126) & x(132) & x(136) & x(152) & x(154) & x(162) & x(180) & x(187) & x(194) & x(207) & x(216) & x(230) & x(236) & x(239) & x(243) & x(244);
    y(42) <= not(p42_out);
    p42 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100001010111011010010010111",
            TABLE => "1000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010010000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010011101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010010001011100000001000101111000000110010110011010010000000000000000",
            SHIFT => 3,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p42_in,
            y(0) => p42_out,
            y(1 to 13 - 1) => dummy42
        );


    p43_in <= x(7) & x(14) & x(16) & x(30) & x(47) & x(51) & x(58) & x(59) & x(72) & x(77) & x(89) & x(90) & x(100) & x(101) & x(123) & x(124) & x(127) & x(130) & x(134) & x(143) & x(212) & x(213) & x(218) & x(224) & x(234) & x(248) & x(254);
    y(43) <= not(p43_out);
    p43 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100011010000100110001101010",
            TABLE => "011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p43_in,
            y(0) => p43_out,
            y(1 to 14 - 1) => dummy43
        );


    p44_in <= x(1) & x(4) & x(5) & x(12) & x(14) & x(17) & x(22) & x(44) & x(52) & x(56) & x(62) & x(66) & x(71) & x(76) & x(85) & x(92) & x(99) & x(100) & x(112) & x(122) & x(123) & x(124) & x(125) & x(142) & x(162) & x(170) & x(174) & x(177) & x(182) & x(206) & x(209) & x(211) & x(217) & x(236) & x(245) & x(247);
    y(44) <= not(p44_out);
    p44 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000101100100010101000110010000110100",
            TABLE => "110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p44_in,
            y(0) => p44_out,
            y(1 to 14 - 1) => dummy44
        );


    p45_in <= x(27) & x(34) & x(39) & x(52) & x(61) & x(62) & x(67) & x(71) & x(77) & x(99) & x(100) & x(102) & x(119) & x(122) & x(123) & x(125) & x(130) & x(144) & x(171) & x(176) & x(182) & x(186) & x(241);
    y(45) <= not(p45_out);
    p45 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00100000100000101111010",
            TABLE => "11101000111111101000000011101000100000001110100000000000100000001110100001111110100000011110100010000001111010000001011110000001011010011001011010010110011010011001011001101001011010011001011011101000111111101000000011101000100000001110100000000000100000001110100001111110100000011110100010000001111010000001011110000001011010011001011010010110011010011001011001101001011010011001011001110001111101110001000001110001000100000111000100000000000100000111000111100111000110000111000100011000011100011000111000011000011010011001011010010110011010011001011001101001011010011001011000100000101100101011001011111011001001001011001010110010110110110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p45_in,
            y(0) => p45_out,
            y(1 to 14 - 1) => dummy45
        );


    p46_in <= x(11) & x(34) & x(57) & x(84) & x(87) & x(93) & x(121) & x(144) & x(148) & x(177) & x(182) & x(215) & x(218);
    y(46) <= not(p46_out);
    p46 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000101100011",
            TABLE => "1111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p46_in,
            y(0) => p46_out,
            y(1 to 13 - 1) => dummy46
        );


    p47_in <= x(11) & x(22) & x(44) & x(56) & x(70) & x(83) & x(89) & x(91) & x(103) & x(135) & x(171) & x(180) & x(183) & x(193) & x(247);
    y(47) <= not(p47_out);
    p47 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010101010101110",
            TABLE => "010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110001010110110100111111111",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p47_in,
            y(0) => p47_out,
            y(1 to 13 - 1) => dummy47
        );


    p48_in <= x(12) & x(17) & x(39) & x(46) & x(63) & x(70) & x(85) & x(102) & x(108) & x(111) & x(114) & x(139) & x(143) & x(153) & x(156) & x(166) & x(178) & x(179) & x(184) & x(187) & x(196) & x(201) & x(202) & x(205) & x(233) & x(236) & x(251);
    y(48) <= not(p48_out);
    p48 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011010100011100100001011101",
            TABLE => "001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110010011010110100111111111",
            SHIFT => 3,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p48_in,
            y(0) => p48_out,
            y(1 to 13 - 1) => dummy48
        );


    p49_in <= x(9) & x(12) & x(22) & x(33) & x(35) & x(48) & x(60) & x(64) & x(75) & x(81) & x(89) & x(101) & x(108) & x(112) & x(123) & x(135) & x(149) & x(151) & x(156) & x(164) & x(178) & x(183) & x(206) & x(231) & x(232) & x(254);
    y(49) <= not(p49_out);
    p49 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00111110110100010001010010",
            TABLE => "000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 3,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p49_in,
            y(0) => p49_out,
            y(1 to 13 - 1) => dummy49
        );


    p50_in <= x(3) & x(4) & x(10) & x(18) & x(25) & x(37) & x(51) & x(53) & x(54) & x(56) & x(58) & x(68) & x(72) & x(76) & x(77) & x(99) & x(101) & x(115) & x(128) & x(131) & x(154) & x(156) & x(160) & x(162) & x(163) & x(171) & x(177) & x(180) & x(182) & x(186) & x(188) & x(189) & x(191) & x(194) & x(206) & x(207);
    y(50) <= not(p50_out);
    p50 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110001110000100111100101101010001110",
            TABLE => "010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p50_in,
            y(0) => p50_out,
            y(1 to 14 - 1) => dummy50
        );


    p51_in <= x(2) & x(26) & x(44) & x(45) & x(64) & x(67) & x(69) & x(73) & x(81) & x(83) & x(90) & x(103) & x(104) & x(120) & x(126) & x(128) & x(157) & x(167) & x(171) & x(174) & x(183) & x(196) & x(201) & x(212) & x(243) & x(252);
    y(51) <= not(p51_out);
    p51 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10100001100101001010010100",
            TABLE => "100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 3,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p51_in,
            y(0) => p51_out,
            y(1 to 13 - 1) => dummy51
        );


    p52_in <= x(3) & x(9) & x(12) & x(33) & x(34) & x(36) & x(50) & x(62) & x(82) & x(86) & x(97) & x(113) & x(115) & x(129) & x(131) & x(134) & x(141) & x(146) & x(163) & x(165) & x(172) & x(188) & x(191) & x(199) & x(205) & x(212) & x(213) & x(216);
    y(52) <= not(p52_out);
    p52 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000110101000010010011001101",
            TABLE => "1111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010011000111000001000111011111000111000001000000000001000111000001000100011100001100011100111100011100001100001110001100011100001100010010110011010010110100110010110011010011001011010010110011010011101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010011000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010000010001001101001001000100110110010110011010010000000000000000",
            SHIFT => 3,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p52_in,
            y(0) => p52_out,
            y(1 to 13 - 1) => dummy52
        );


    p53_in <= x(3) & x(4) & x(35) & x(36) & x(58) & x(82) & x(126) & x(130) & x(132) & x(133) & x(134) & x(158) & x(160) & x(163) & x(171) & x(181) & x(189) & x(203) & x(208) & x(211) & x(227) & x(230) & x(243) & x(244);
    y(53) <= not(p53_out);
    p53 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100111100011110100010111",
            TABLE => "000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p53_in,
            y(0) => p53_out,
            y(1 to 14 - 1) => dummy53
        );


    p54_in <= x(5) & x(26) & x(48) & x(67) & x(70) & x(79) & x(87) & x(101) & x(106) & x(123) & x(127) & x(129) & x(130) & x(133) & x(140) & x(149) & x(174) & x(198) & x(205) & x(217) & x(218) & x(230) & x(254);
    y(54) <= not(p54_out);
    p54 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11110011101011001111000",
            TABLE => "00000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100100000000001000000010000010110010001000001011001010110010111110110100110100100100001001001011001000100100101100101011001011011011100101100110100101101001100101100110100110010110100101100110100100010000000000000111000100010000011100010001000011110111011100010001100010001110011100010001100001110001000110001110011101110001100101100110100101101001100101100110100110010110100101100110100110000000111010001110100011111110100000011110100011101000011111101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p54_in,
            y(0) => p54_out,
            y(1 to 14 - 1) => dummy54
        );


    p55_in <= x(4) & x(15) & x(21) & x(36) & x(47) & x(52) & x(95) & x(103) & x(108) & x(110) & x(114) & x(129) & x(134) & x(140) & x(141) & x(143) & x(164) & x(165) & x(181) & x(189) & x(197) & x(219) & x(224) & x(230) & x(235) & x(236) & x(238) & x(243) & x(247);
    y(55) <= not(p55_out);
    p55 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00110101001000011000110011000",
            TABLE => "01001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011010110010001000001111101110110010001000000000000010110010001000001011001000100100110110111011001000100100010011011011001000100100100101100110100101101001100101100110100110010110100101100110100110111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100110001110111011110000100010001110000010001000111000000000000010001000111011100111000110001000111000011000100011100111000100011000100101100110100101101001100101100110100110010110100101100110100110000000111010001110100011111110100000011110100011101000011111101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p55_in,
            y(0) => p55_out,
            y(1 to 14 - 1) => dummy55
        );


    p56_in <= x(4) & x(33) & x(51) & x(55) & x(56) & x(57) & x(60) & x(70) & x(79) & x(80) & x(83) & x(86) & x(89) & x(91) & x(99) & x(101) & x(117) & x(123) & x(129) & x(131) & x(133) & x(140) & x(151) & x(166) & x(172) & x(179) & x(182) & x(194) & x(199) & x(218) & x(238) & x(246) & x(248) & x(253) & x(255);
    y(56) <= not(p56_out);
    p56 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10010101100110001101011010100111001",
            TABLE => "01001101000001000000010000000000110111110100110101001101000001000100110100100100001001001011001011011011010011010100110100100100011010011001011010010110011010011001011001101001011010011001011001000000110101001101010011111101000000000100000001000000110101000100001011010100110101001011110100101011010000100100001011010100011010011001011010010110011010011001011001101001011010011001011001110001000100000001000000000000111101110111000101110001000100000111000100011000000110001000111011100111011100010111000100011000011010011001011010010110011010011001011001101001011010011001011000101011000000101011111100101011000000100000000000101011000000100010101101000010101111010010101101000010110101000010101101000010011010011001011010010110011010011001011001101001011010011001011001000000110101000000000001000000110101001111110101000000110101000100001011010100001010110100001011010100101111010100001011010100011010011001011010010110011010011001011001101001011010011001011001000000110101001101010011111101010000101101010011010100101111010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 3,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p56_in,
            y(0) => p56_out,
            y(1 to 14 - 1) => dummy56
        );


    p57_in <= x(12) & x(35) & x(36) & x(47) & x(71) & x(79) & x(85) & x(92) & x(93) & x(103) & x(105) & x(114) & x(119) & x(143) & x(151) & x(160) & x(168) & x(177) & x(180) & x(182) & x(186) & x(190) & x(202) & x(207) & x(219) & x(231) & x(237) & x(240);
    y(57) <= not(p57_out);
    p57 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101010100000011001011010111",
            TABLE => "0000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010011110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101101000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010001011100000001000101111000000110010110011010010000000000000000",
            SHIFT => 3,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p57_in,
            y(0) => p57_out,
            y(1 to 13 - 1) => dummy57
        );


    p58_in <= x(4) & x(15) & x(26) & x(51) & x(56) & x(58) & x(86) & x(89) & x(94) & x(101) & x(106) & x(118) & x(129) & x(131) & x(145) & x(156) & x(166) & x(170) & x(179) & x(191) & x(192) & x(203) & x(213) & x(215) & x(218) & x(246) & x(248) & x(252);
    y(58) <= not(p58_out);
    p58 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001100001111011101111100010",
            TABLE => "1011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101011001000100000101100100010010010010110011010010000000000000000",
            SHIFT => 3,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p58_in,
            y(0) => p58_out,
            y(1 to 13 - 1) => dummy58
        );


    p59_in <= x(5) & x(15) & x(31) & x(48) & x(56) & x(57) & x(60) & x(66) & x(80) & x(87) & x(89) & x(94) & x(102) & x(131) & x(139) & x(140) & x(149) & x(151) & x(162) & x(166) & x(168) & x(176) & x(179) & x(192) & x(195) & x(212) & x(234) & x(236) & x(241) & x(244) & x(248) & x(249);
    y(59) <= not(p59_out);
    p59 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01000101001111011100100010111001",
            TABLE => "110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p59_in,
            y(0) => p59_out,
            y(1 to 14 - 1) => dummy59
        );


    p60_in <= x(4) & x(6) & x(24) & x(26) & x(47) & x(56) & x(62) & x(76) & x(77) & x(93) & x(99) & x(119) & x(122) & x(129) & x(135) & x(140) & x(149) & x(151) & x(160) & x(164) & x(169) & x(173) & x(180) & x(182) & x(183) & x(202) & x(207) & x(214) & x(219) & x(223) & x(224) & x(240) & x(248) & x(254);
    y(60) <= not(p60_out);
    p60 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001001001111010000111011100101000",
            TABLE => "1000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010011000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101101000000011101000100000011110100010010110011010010000000000000000",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p60_in,
            y(0) => p60_out,
            y(1 to 14 - 1) => dummy60
        );


    p61_in <= x(3) & x(4) & x(14) & x(45) & x(85) & x(87) & x(105) & x(110) & x(114) & x(129) & x(152) & x(153) & x(157) & x(158) & x(159) & x(160) & x(181) & x(202) & x(208) & x(211) & x(223) & x(226) & x(235) & x(236) & x(248);
    y(61) <= not(p61_out);
    p61 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111010000100001001011101",
            TABLE => "0000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101101110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p61_in,
            y(0) => p61_out,
            y(1 to 14 - 1) => dummy61
        );


    p62_in <= x(9) & x(18) & x(19) & x(21) & x(26) & x(29) & x(37) & x(50) & x(58) & x(63) & x(75) & x(81) & x(89) & x(101) & x(102) & x(113) & x(131) & x(138) & x(140) & x(141) & x(160) & x(163) & x(179) & x(181) & x(188) & x(191) & x(192) & x(195) & x(196) & x(207) & x(213) & x(234) & x(236) & x(239);
    y(62) <= not(p62_out);
    p62 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111110010111010111010011001010100",
            TABLE => "0000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101100001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010010100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101101000111000001000100011100001100010010110011010010000000000000000",
            SHIFT => 3,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p62_in,
            y(0) => p62_out,
            y(1 to 14 - 1) => dummy62
        );


    p63_in <= x(10) & x(15) & x(21) & x(40) & x(44) & x(48) & x(59) & x(61) & x(78) & x(80) & x(86) & x(89) & x(90) & x(127) & x(133) & x(135) & x(138) & x(139) & x(145) & x(148) & x(151) & x(156) & x(161) & x(162) & x(164) & x(167) & x(177) & x(183) & x(185) & x(190) & x(203) & x(205) & x(209) & x(210) & x(216) & x(223) & x(235) & x(245) & x(248) & x(255);
    y(63) <= not(p63_out);
    p63 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000101011001010011011010010101000111110",
            TABLE => "1111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100000100010001110000000000000100010001110111011110000100010001110000110001000111001110001000110001000111011100111000110001000111001101001100101101001011001101001100101100110100101101001100101100100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010011011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010010111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101100000001000101011010000100010101110010110011010010000000000000000",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p63_in,
            y(0) => p63_out,
            y(1 to 15 - 1) => dummy63
        );


    p64_in <= x(18) & x(34) & x(39) & x(55) & x(78) & x(81) & x(99) & x(100) & x(101) & x(102) & x(103) & x(107) & x(113) & x(131) & x(148) & x(152) & x(160) & x(168) & x(173) & x(174) & x(184) & x(186) & x(190) & x(200) & x(203) & x(204) & x(209) & x(219) & x(224) & x(232) & x(237) & x(241) & x(242);
    y(64) <= not(p64_out);
    p64 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010000111111001101111000000111010",
            TABLE => "111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => 3,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p64_in,
            y(0) => p64_out,
            y(1 to 14 - 1) => dummy64
        );


    p65_in <= x(1) & x(3) & x(4) & x(11) & x(13) & x(14) & x(18) & x(29) & x(37) & x(38) & x(45) & x(46) & x(49) & x(88) & x(95) & x(98) & x(104) & x(110) & x(112) & x(130) & x(137) & x(140) & x(144) & x(175) & x(196) & x(207) & x(208) & x(209) & x(214) & x(216) & x(229) & x(230) & x(236) & x(250) & x(251) & x(255);
    y(65) <= not(p65_out);
    p65 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011000101101110100011010101001001110",
            TABLE => "100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p65_in,
            y(0) => p65_out,
            y(1 to 14 - 1) => dummy65
        );


    p66_in <= x(4) & x(10) & x(28) & x(29) & x(63) & x(64) & x(79) & x(81) & x(108) & x(173) & x(178) & x(196) & x(201) & x(213) & x(224);
    y(66) <= not(p66_out);
    p66 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010010010001000",
            TABLE => "101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p66_in,
            y(0) => p66_out,
            y(1 to 13 - 1) => dummy66
        );


    p67_in <= x(3) & x(9) & x(28) & x(30) & x(34) & x(37) & x(49) & x(50) & x(77) & x(78) & x(94) & x(103) & x(104) & x(111) & x(120) & x(134) & x(146) & x(149) & x(155) & x(188) & x(199) & x(212) & x(222) & x(224) & x(232) & x(233) & x(254);
    y(67) <= not(p67_out);
    p67 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001010000001111010110101100",
            TABLE => "101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001100011101001011011111111",
            SHIFT => 3,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p67_in,
            y(0) => p67_out,
            y(1 to 13 - 1) => dummy67
        );


    p68_in <= x(33) & x(53) & x(71) & x(72) & x(74) & x(77) & x(83) & x(103) & x(105) & x(120) & x(123) & x(165) & x(168) & x(174) & x(179) & x(188) & x(194) & x(199) & x(209) & x(212) & x(252) & x(253) & x(254);
    y(68) <= not(p68_out);
    p68 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001001111000110011000",
            TABLE => "11111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011000000010001010110010101110111111000000000000001000000010001010110100001000101011001010111011110111010100010000100100001000101011100101100110100101101001100101100110100110010110100101100110100110001110111011110000100010001110000010001000111000000000000010001000111011100111000110001000111000011000100011100111000100011000100101100110100101101001100101100110100110010110100101100110100110000000111010001110100011111110100000011110100011101000011111101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p68_in,
            y(0) => p68_out,
            y(1 to 14 - 1) => dummy68
        );


    p69_in <= x(4) & x(6) & x(7) & x(8) & x(17) & x(19) & x(28) & x(53) & x(96) & x(104) & x(135) & x(147) & x(153) & x(163) & x(164) & x(173) & x(183) & x(193) & x(214) & x(219) & x(235) & x(254);
    y(69) <= not(p69_out);
    p69 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111000110011100001001",
            TABLE => "0000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101101000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010100000011010100010000101101010001101001100101100000000000000000",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p69_in,
            y(0) => p69_out,
            y(1 to 14 - 1) => dummy69
        );


    p70_in <= x(9) & x(10) & x(17) & x(22) & x(24) & x(32) & x(58) & x(74) & x(77) & x(99) & x(109) & x(131) & x(139) & x(141) & x(150) & x(155) & x(163) & x(168) & x(171) & x(176) & x(191) & x(199) & x(203) & x(206) & x(207) & x(213) & x(225) & x(230) & x(239);
    y(70) <= not(p70_out);
    p70 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10010000010011101100110101111",
            TABLE => "10001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100111101111100011101000111000001000100011100000100000001000000000001110011110001110100011100001100010001110000110000001100001110001011010011001011010010110011010011001011001101001011010011001011000000000000100000001000001110001000100000111000101110001111101111000111000011000000110000111000100011000011100010111000111100111011010011001011010010110011010011001011001101001011010011001011001001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011000010111011111110000000100010111000101110111111010000001000101111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p70_in,
            y(0) => p70_out,
            y(1 to 14 - 1) => dummy70
        );


    p71_in <= x(5) & x(7) & x(25) & x(32) & x(35) & x(39) & x(53) & x(62) & x(63) & x(64) & x(69) & x(82) & x(89) & x(91) & x(99) & x(100) & x(102) & x(137) & x(143) & x(149) & x(150) & x(158) & x(161) & x(162) & x(183) & x(184) & x(193) & x(197) & x(207) & x(216) & x(232) & x(234) & x(245);
    y(71) <= not(p71_out);
    p71 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110100111000101000111001000101001",
            TABLE => "000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001110101001001011011111111",
            SHIFT => 4,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p71_in,
            y(0) => p71_out,
            y(1 to 15 - 1) => dummy71
        );


    p72_in <= x(4) & x(12) & x(17) & x(25) & x(38) & x(42) & x(46) & x(47) & x(82) & x(98) & x(111) & x(115) & x(118) & x(135) & x(139) & x(151) & x(153) & x(158) & x(177) & x(187) & x(192) & x(196) & x(219) & x(221) & x(224) & x(227) & x(232) & x(234) & x(235) & x(236) & x(251);
    y(72) <= not(p72_out);
    p72 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100001101101001101100011100010",
            TABLE => "1000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010010010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101100100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p72_in,
            y(0) => p72_out,
            y(1 to 14 - 1) => dummy72
        );


    p73_in <= x(5) & x(16) & x(29) & x(39) & x(40) & x(59) & x(68) & x(72) & x(74) & x(80) & x(86) & x(117) & x(129) & x(137) & x(162) & x(227) & x(230) & x(244) & x(247) & x(249);
    y(73) <= not(p73_out);
    p73 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01001010101101010001",
            TABLE => "101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 4,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p73_in,
            y(0) => p73_out,
            y(1 to 14 - 1) => dummy73
        );


    p74_in <= x(4) & x(14) & x(34) & x(40) & x(44) & x(50) & x(55) & x(56) & x(62) & x(65) & x(67) & x(74) & x(79) & x(90) & x(91) & x(104) & x(113) & x(123) & x(126) & x(129) & x(139) & x(156) & x(160) & x(167) & x(168) & x(171) & x(179) & x(186) & x(204) & x(205) & x(212) & x(218) & x(231) & x(253);
    y(74) <= not(p74_out);
    p74 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0011000101110111001101111010000001",
            TABLE => "1000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010010000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101101000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010011101010001000000110101000100001010010110011010010000000000000000",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p74_in,
            y(0) => p74_out,
            y(1 to 15 - 1) => dummy74
        );


    p75_in <= x(5) & x(26) & x(52) & x(79) & x(95) & x(108) & x(119) & x(125) & x(126) & x(130) & x(134) & x(136) & x(141) & x(154) & x(160) & x(163) & x(178) & x(182) & x(184) & x(191) & x(197) & x(214) & x(218) & x(220) & x(232) & x(235) & x(236) & x(238) & x(241) & x(243) & x(246) & x(253);
    y(75) <= not(p75_out);
    p75 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00011101101110111111011010111110",
            TABLE => "011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p75_in,
            y(0) => p75_out,
            y(1 to 14 - 1) => dummy75
        );


    p76_in <= x(4) & x(7) & x(8) & x(12) & x(16) & x(51) & x(64) & x(73) & x(81) & x(87) & x(108) & x(118) & x(129) & x(133) & x(151) & x(158) & x(159) & x(170) & x(182) & x(193) & x(197) & x(211) & x(217) & x(226) & x(235) & x(240) & x(246) & x(248);
    y(76) <= not(p76_out);
    p76 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110010111010110000010111101",
            TABLE => "0100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010011000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101100000010001001101001001000100110110010110011010010000000000000000",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p76_in,
            y(0) => p76_out,
            y(1 to 13 - 1) => dummy76
        );


    p77_in <= x(3) & x(25) & x(33) & x(37) & x(59) & x(60) & x(93) & x(101) & x(104) & x(115) & x(121) & x(131) & x(146) & x(159) & x(163) & x(168) & x(174) & x(203) & x(206) & x(212) & x(223) & x(226) & x(235) & x(240) & x(241) & x(242) & x(252);
    y(77) <= not(p77_out);
    p77 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101100011110011110100000101",
            TABLE => "000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110010011010110100111111111",
            SHIFT => 3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p77_in,
            y(0) => p77_out,
            y(1 to 13 - 1) => dummy77
        );


    p78_in <= x(16) & x(26) & x(29) & x(33) & x(34) & x(37) & x(65) & x(75) & x(78) & x(100) & x(130) & x(154) & x(165) & x(167) & x(168) & x(181) & x(184) & x(197) & x(198) & x(200) & x(212) & x(232) & x(240) & x(243) & x(250) & x(253);
    y(78) <= not(p78_out);
    p78 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01010110101111100111000011",
            TABLE => "010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p78_in,
            y(0) => p78_out,
            y(1 to 14 - 1) => dummy78
        );


    p79_in <= x(9) & x(18) & x(37) & x(52) & x(59) & x(62) & x(67) & x(88) & x(115) & x(125) & x(139) & x(147) & x(151) & x(160) & x(165) & x(173) & x(200) & x(236);
    y(79) <= not(p79_out);
    p79 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101001111110001110",
            TABLE => "010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p79_in,
            y(0) => p79_out,
            y(1 to 14 - 1) => dummy79
        );


    p80_in <= x(5) & x(12) & x(32) & x(39) & x(41) & x(46) & x(48) & x(62) & x(64) & x(70) & x(77) & x(87) & x(94) & x(108) & x(113) & x(115) & x(117) & x(119) & x(120) & x(130) & x(136) & x(137) & x(147) & x(149) & x(151) & x(153) & x(162) & x(190) & x(194) & x(236) & x(242) & x(249);
    y(80) <= not(p80_out);
    p80 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01001100110011001000011111010101",
            TABLE => "011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 3,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p80_in,
            y(0) => p80_out,
            y(1 to 14 - 1) => dummy80
        );


    p81_in <= x(7) & x(14) & x(25) & x(39) & x(42) & x(44) & x(47) & x(50) & x(51) & x(98) & x(114) & x(115) & x(118) & x(119) & x(140) & x(143) & x(151) & x(158) & x(164) & x(166) & x(211) & x(227) & x(232) & x(247);
    y(81) <= not(p81_out);
    p81 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110001101100101010000101",
            TABLE => "010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p81_in,
            y(0) => p81_out,
            y(1 to 14 - 1) => dummy81
        );


    p82_in <= x(9) & x(10) & x(11) & x(18) & x(24) & x(44) & x(49) & x(52) & x(55) & x(61) & x(63) & x(65) & x(66) & x(67) & x(69) & x(73) & x(74) & x(77) & x(81) & x(99) & x(105) & x(125) & x(128) & x(145) & x(160) & x(165) & x(167) & x(173) & x(175) & x(183) & x(187) & x(213) & x(222) & x(239) & x(249);
    y(82) <= not(p82_out);
    p82 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01111100100000011110100110001010001",
            TABLE => "00000001000101110001011101111111000000000000000100000001000101111000000100010111000101110111111011101000100000011000000100010111011010011001011010010110011010011001011001101001011010011001011011101000111111101000000011101000100000001110100000000000100000001110100001111110100000011110100010000001111010000001011110000001011010011001011010010110011010011001011001101001011010011001011001111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011001000000110101000000000001000000110101001111110101000000110101000100001011010100001010110100001011010100101111010100001011010100011010011001011010010110011010011001011001101001011010011001011010110010001000000010000000000000111110111011001010110010001000001011001000100100001001000100110111011011101100101011001000100100100101100110100101101001100101100110100110010110100101100110100111010100010000001111110111010100110101000100001010111101110101001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p82_in,
            y(0) => p82_out,
            y(1 to 14 - 1) => dummy82
        );


    p83_in <= x(1) & x(3) & x(4) & x(12) & x(40) & x(49) & x(52) & x(53) & x(71) & x(72) & x(79) & x(92) & x(106) & x(108) & x(114) & x(119) & x(122) & x(130) & x(166) & x(168) & x(176) & x(178) & x(186) & x(204) & x(226) & x(235) & x(242);
    y(83) <= not(p83_out);
    p83 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001100000011010001001111111",
            TABLE => "100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 3,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p83_in,
            y(0) => p83_out,
            y(1 to 13 - 1) => dummy83
        );


    p84_in <= x(18) & x(20) & x(26) & x(28) & x(44) & x(48) & x(66) & x(67) & x(68) & x(87) & x(94) & x(95) & x(101) & x(110) & x(129) & x(133) & x(136) & x(154) & x(162) & x(163) & x(175) & x(180) & x(181) & x(191) & x(195) & x(207) & x(208) & x(215) & x(226) & x(230) & x(234) & x(243) & x(247) & x(253);
    y(84) <= not(p84_out);
    p84 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0101110000011110101110110000010110",
            TABLE => "0001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010010000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101101111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p84_in,
            y(0) => p84_out,
            y(1 to 14 - 1) => dummy84
        );


    p85_in <= x(15) & x(23) & x(28) & x(32) & x(40) & x(49) & x(55) & x(68) & x(113) & x(137) & x(162) & x(168) & x(172) & x(175) & x(176) & x(180) & x(181) & x(195) & x(200) & x(202) & x(204) & x(209) & x(227) & x(244);
    y(85) <= not(p85_out);
    p85 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001100101010111010111101",
            TABLE => "100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p85_in,
            y(0) => p85_out,
            y(1 to 13 - 1) => dummy85
        );


    p86_in <= x(12) & x(20) & x(26) & x(28) & x(30) & x(34) & x(37) & x(44) & x(48) & x(70) & x(73) & x(94) & x(103) & x(105) & x(120) & x(146) & x(150) & x(181) & x(182) & x(199) & x(201);
    y(86) <= not(p86_out);
    p86 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101010100101000010011",
            TABLE => "001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p86_in,
            y(0) => p86_out,
            y(1 to 14 - 1) => dummy86
        );


    p87_in <= x(3) & x(10) & x(32) & x(35) & x(37) & x(60) & x(61) & x(71) & x(83) & x(95) & x(103) & x(116) & x(126) & x(160) & x(182) & x(202) & x(206) & x(207) & x(216) & x(223) & x(225) & x(237) & x(240);
    y(87) <= not(p87_out);
    p87 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110100110111000101011",
            TABLE => "00000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100101001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011001000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011001110001111101110001000001110001011100011110011100011000011100010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p87_in,
            y(0) => p87_out,
            y(1 to 14 - 1) => dummy87
        );


    p88_in <= x(22) & x(32) & x(37) & x(39) & x(42) & x(46) & x(47) & x(51) & x(54) & x(60) & x(82) & x(90) & x(95) & x(96) & x(98) & x(112) & x(113) & x(118) & x(121) & x(134) & x(151) & x(172) & x(174) & x(175) & x(195) & x(203) & x(204) & x(209) & x(216) & x(222) & x(228) & x(231) & x(234) & x(237) & x(241) & x(242) & x(248);
    y(88) <= not(p88_out);
    p88 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010011100000110011010101000100000101",
            TABLE => "0100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101101000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101101011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 3,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p88_in,
            y(0) => p88_out,
            y(1 to 14 - 1) => dummy88
        );


    p89_in <= x(9) & x(23) & x(25) & x(26) & x(52) & x(55) & x(56) & x(66) & x(82) & x(89) & x(92) & x(93) & x(94) & x(96) & x(107) & x(122) & x(128) & x(129) & x(131) & x(139) & x(157) & x(186) & x(191) & x(192) & x(197) & x(199) & x(201) & x(211) & x(213) & x(220) & x(225) & x(228) & x(232) & x(234) & x(242) & x(245) & x(252);
    y(89) <= not(p89_out);
    p89 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010011010100110010111110001101110100",
            TABLE => "0100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101100100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101101011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010010000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p89_in,
            y(0) => p89_out,
            y(1 to 14 - 1) => dummy89
        );


    p90_in <= x(9) & x(12) & x(13) & x(28) & x(37) & x(38) & x(49) & x(52) & x(65) & x(66) & x(79) & x(82) & x(93) & x(95) & x(103) & x(110) & x(112) & x(113) & x(143) & x(161) & x(162) & x(163) & x(168) & x(173) & x(178) & x(192) & x(193) & x(197) & x(216) & x(237) & x(243) & x(253);
    y(90) <= not(p90_out);
    p90 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001111110010100011001000011001",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 3,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p90_in,
            y(0) => p90_out,
            y(1 to 14 - 1) => dummy90
        );


    p91_in <= x(12) & x(35) & x(37) & x(40) & x(45) & x(52) & x(54) & x(62) & x(63) & x(65) & x(66) & x(76) & x(78) & x(93) & x(100) & x(102) & x(103) & x(124) & x(133) & x(140) & x(142) & x(160) & x(162) & x(183) & x(184) & x(193) & x(196) & x(197) & x(216) & x(232) & x(234) & x(247) & x(249) & x(250) & x(251);
    y(91) <= not(p91_out);
    p91 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11011010000100110101010111000110100",
            TABLE => "00000010000000000010101100000010001010110000001010111111001010110100001011010100001010110100001000101011010000101011110100101011100101100110100101101001100101100110100110010110100101100110100111010100010000000100000000000000111111011101010011010100010000001101010001000010010000100010101110111101110101001101010001000010100101100110100101101001100101100110100110010110100101100110100101001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011001001101000001001101111101001101000001000000000001001101000001000100110100100100110110110100110100100100101100100100110100100100011010011001011010010110011010011001011001101001011010011001011001000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011010001110000010001110111110001110100011100001100011100111100011101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p91_in,
            y(0) => p91_out,
            y(1 to 15 - 1) => dummy91
        );


    p92_in <= x(14) & x(28) & x(31) & x(40) & x(41) & x(47) & x(62) & x(72) & x(90) & x(98) & x(103) & x(119) & x(121) & x(132) & x(139) & x(142) & x(152) & x(169) & x(205) & x(225) & x(227) & x(236) & x(251);
    y(92) <= not(p92_out);
    p92 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11100011101100110010001",
            TABLE => "00000000100000001000000011101000100000001110100011101000111111100001011110000001100000011110100010000001111010001110100001111110011010011001011010010110011010011001011001101001011010011001011000000000000100000001000001110001000100000111000101110001111101111000111000011000000110000111000100011000011100010111000111100111011010011001011010010110011010011001011001101001011010011001011010001110111011110000100010001110000010001000111000000000000010001000111011100111000110001000111000011000100011100111000100011000100101100110100101101001100101100110100110010110100101100110100111010100010000001111110111010100110101000100001010111101110101001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p92_in,
            y(0) => p92_out,
            y(1 to 14 - 1) => dummy92
        );


    p93_in <= x(2) & x(14) & x(26) & x(40) & x(50) & x(59) & x(63) & x(67) & x(79) & x(80) & x(112) & x(134) & x(136) & x(137) & x(154) & x(172) & x(176) & x(189) & x(195) & x(224) & x(248) & x(253);
    y(93) <= not(p93_out);
    p93 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1011010101000010001011",
            TABLE => "0000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010011000111000001000111011111000111000001000000000001000111000001000100011100001100011100111100011100001100001110001100011100001100010010110011010010110100110010110011010011001011010010110011010011110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100001000001110001000110000111000110010110011010010000000000000000",
            SHIFT => 4,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p93_in,
            y(0) => p93_out,
            y(1 to 14 - 1) => dummy93
        );


    p94_in <= x(0) & x(1) & x(8) & x(10) & x(14) & x(28) & x(44) & x(72) & x(75) & x(88) & x(89) & x(93) & x(95) & x(108) & x(109) & x(111) & x(136) & x(137) & x(145) & x(147) & x(156) & x(157) & x(160) & x(164) & x(166) & x(180) & x(184) & x(197) & x(211) & x(214) & x(224) & x(232) & x(235) & x(238) & x(241) & x(254) & x(255);
    y(94) <= not(p94_out);
    p94 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111101110101010101100101001010001111",
            TABLE => "0000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010010010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101100010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101100100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 3,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p94_in,
            y(0) => p94_out,
            y(1 to 14 - 1) => dummy94
        );


    p95_in <= x(14) & x(22) & x(26) & x(36) & x(44) & x(59) & x(61) & x(64) & x(67) & x(76) & x(112) & x(127) & x(136) & x(142) & x(145) & x(149) & x(154) & x(164) & x(173) & x(198) & x(226) & x(231) & x(254);
    y(95) <= not(p95_out);
    p95 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10011001001011110010011",
            TABLE => "00101011000000100000001000000000101111110010101100101011000000100010101101000010010000101101010010111101001010110010101101000010011010011001011010010110011010011001011001101001011010011001011010110010001000001111101110110010001000000000000010110010001000001011001000100100110110111011001000100100010011011011001000100100100101100110100101101001100101100110100110010110100101100110100100000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100101110001000100001111011101110001011100010001100011100111011100010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p95_in,
            y(0) => p95_out,
            y(1 to 14 - 1) => dummy95
        );


    p96_in <= x(2) & x(7) & x(8) & x(10) & x(18) & x(27) & x(29) & x(52) & x(64) & x(67) & x(69) & x(73) & x(78) & x(81) & x(88) & x(100) & x(102) & x(124) & x(126) & x(130) & x(144) & x(148) & x(156) & x(166) & x(171) & x(178) & x(182) & x(183) & x(184) & x(220) & x(232) & x(243) & x(248);
    y(96) <= not(p96_out);
    p96 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000001101110001110100110011110110",
            TABLE => "111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001001010110110100111111111",
            SHIFT => 3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p96_in,
            y(0) => p96_out,
            y(1 to 14 - 1) => dummy96
        );


    p97_in <= x(27) & x(28) & x(34) & x(49) & x(77) & x(78) & x(87) & x(107) & x(111) & x(120) & x(121) & x(127) & x(130) & x(142) & x(148) & x(153) & x(179) & x(183) & x(184) & x(188) & x(199) & x(212) & x(220) & x(222) & x(231) & x(232) & x(242) & x(246);
    y(97) <= not(p97_out);
    p97 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001111000101100000010111010",
            TABLE => "0111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101101011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010011000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101100010000010110010001001001011001001101001100101100000000000000000",
            SHIFT => 3,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p97_in,
            y(0) => p97_out,
            y(1 to 13 - 1) => dummy97
        );


    p98_in <= x(1) & x(3) & x(4) & x(6) & x(7) & x(11) & x(26) & x(38) & x(45) & x(47) & x(63) & x(65) & x(76) & x(89) & x(91) & x(107) & x(114) & x(118) & x(119) & x(132) & x(135) & x(139) & x(140) & x(142) & x(150) & x(157) & x(158) & x(162) & x(166) & x(174) & x(192) & x(196) & x(224) & x(227) & x(228) & x(229) & x(232) & x(241);
    y(98) <= not(p98_out);
    p98 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10101110110101000101001110010100110101",
            TABLE => "000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 3,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p98_in,
            y(0) => p98_out,
            y(1 to 14 - 1) => dummy98
        );


    p99_in <= x(14) & x(39) & x(40) & x(55) & x(56) & x(59) & x(63) & x(67) & x(83) & x(85) & x(103) & x(109) & x(123) & x(126) & x(127) & x(151) & x(161) & x(180) & x(182) & x(193) & x(206) & x(216) & x(218) & x(225) & x(247);
    y(99) <= not(p99_out);
    p99 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001001001101001001011111",
            TABLE => "1000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101101000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p99_in,
            y(0) => p99_out,
            y(1 to 14 - 1) => dummy99
        );


    p100_in <= x(12) & x(15) & x(39) & x(42) & x(46) & x(52) & x(58) & x(69) & x(70) & x(83) & x(95) & x(96) & x(103) & x(111) & x(112) & x(116) & x(136) & x(142) & x(157) & x(167) & x(179) & x(184) & x(187) & x(191) & x(207) & x(220) & x(225) & x(232) & x(242) & x(252);
    y(100) <= not(p100_out);
    p100 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001101110110001111010000110011",
            TABLE => "010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p100_in,
            y(0) => p100_out,
            y(1 to 14 - 1) => dummy100
        );


    p101_in <= x(8) & x(29) & x(34) & x(37) & x(52) & x(59) & x(63) & x(95) & x(100) & x(104) & x(113) & x(126) & x(150) & x(160) & x(179) & x(184) & x(197) & x(200) & x(205) & x(207) & x(220) & x(228) & x(232) & x(233) & x(240);
    y(101) <= not(p101_out);
    p101 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110010111010111000101101",
            TABLE => "0100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p101_in,
            y(0) => p101_out,
            y(1 to 14 - 1) => dummy101
        );


    p102_in <= x(3) & x(25) & x(36) & x(38) & x(43) & x(47) & x(68) & x(80) & x(87) & x(91) & x(114) & x(115) & x(117) & x(124) & x(128) & x(166) & x(181) & x(186) & x(187) & x(189) & x(206) & x(221) & x(226) & x(230) & x(239) & x(242) & x(249);
    y(102) <= not(p102_out);
    p102 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010001101000110001110110011",
            TABLE => "110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001011100010110100111111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p102_in,
            y(0) => p102_out,
            y(1 to 14 - 1) => dummy102
        );


    p103_in <= x(6) & x(35) & x(47) & x(58) & x(78) & x(115) & x(118) & x(130) & x(132) & x(133) & x(148) & x(158) & x(159) & x(202) & x(213) & x(217) & x(221) & x(232) & x(242) & x(255);
    y(103) <= not(p103_out);
    p103 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10010100001111000101",
            TABLE => "010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p103_in,
            y(0) => p103_out,
            y(1 to 14 - 1) => dummy103
        );


    p104_in <= x(4) & x(5) & x(10) & x(26) & x(33) & x(34) & x(67) & x(74) & x(80) & x(99) & x(107) & x(122) & x(130) & x(132) & x(142) & x(149) & x(161) & x(168) & x(169) & x(188) & x(198) & x(200) & x(224) & x(241) & x(250);
    y(104) <= not(p104_out);
    p104 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010010100100011100100010",
            TABLE => "1101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010011011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010010010101110111111000000100010101100000010001010110000000000000010001010111011110101000010001010110100001000101011110101000100001001101001100101101001011001101001100101100110100101101001100101101101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p104_in,
            y(0) => p104_out,
            y(1 to 14 - 1) => dummy104
        );


    p105_in <= x(1) & x(4) & x(9) & x(11) & x(12) & x(20) & x(43) & x(55) & x(64) & x(76) & x(81) & x(91) & x(92) & x(105) & x(134) & x(141) & x(147) & x(153) & x(178) & x(193) & x(247);
    y(105) <= not(p105_out);
    p105 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011010011101101100110",
            TABLE => "001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110001010110110100111111111",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p105_in,
            y(0) => p105_out,
            y(1 to 14 - 1) => dummy105
        );


    p106_in <= x(0) & x(5) & x(17) & x(28) & x(29) & x(33) & x(40) & x(49) & x(68) & x(75) & x(86) & x(101) & x(103) & x(137) & x(141) & x(166) & x(176) & x(177) & x(182) & x(195) & x(245);
    y(106) <= not(p106_out);
    p106 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001001111010011100010",
            TABLE => "110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => 4,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p106_in,
            y(0) => p106_out,
            y(1 to 14 - 1) => dummy106
        );


    p107_in <= x(25) & x(41) & x(52) & x(53) & x(70) & x(78) & x(82) & x(83) & x(93) & x(100) & x(103) & x(109) & x(110) & x(115) & x(118) & x(126) & x(133) & x(151) & x(158) & x(159) & x(171) & x(181) & x(197) & x(199) & x(216) & x(221) & x(226) & x(235) & x(243) & x(250);
    y(107) <= not(p107_out);
    p107 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000100110101110100110101000010",
            TABLE => "111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p107_in,
            y(0) => p107_out,
            y(1 to 14 - 1) => dummy107
        );


    p108_in <= x(0) & x(1) & x(6) & x(7) & x(19) & x(25) & x(39) & x(78) & x(128) & x(153) & x(157) & x(159) & x(169) & x(180) & x(191) & x(198) & x(204) & x(207) & x(217) & x(225) & x(226) & x(235) & x(240) & x(243);
    y(108) <= not(p108_out);
    p108 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000011110000010011101110",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p108_in,
            y(0) => p108_out,
            y(1 to 14 - 1) => dummy108
        );


    p109_in <= x(0) & x(3) & x(7) & x(15) & x(25) & x(35) & x(53) & x(61) & x(71) & x(72) & x(106) & x(137) & x(139) & x(153) & x(167) & x(175) & x(186) & x(203) & x(206) & x(207) & x(222) & x(223) & x(235) & x(240) & x(242) & x(255);
    y(109) <= not(p109_out);
    p109 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001100000110001101011110",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p109_in,
            y(0) => p109_out,
            y(1 to 14 - 1) => dummy109
        );


    p110_in <= x(5) & x(8) & x(17) & x(25) & x(34) & x(35) & x(63) & x(70) & x(83) & x(103) & x(135) & x(147) & x(149) & x(161) & x(171) & x(186) & x(193) & x(206) & x(207) & x(215) & x(216) & x(228) & x(240) & x(245);
    y(110) <= not(p110_out);
    p110 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110000110101101001001001",
            TABLE => "100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p110_in,
            y(0) => p110_out,
            y(1 to 14 - 1) => dummy110
        );


    p111_in <= x(0) & x(6) & x(12) & x(17) & x(21) & x(26) & x(36) & x(40) & x(44) & x(45) & x(46) & x(47) & x(51) & x(62) & x(77) & x(96) & x(98) & x(103) & x(110) & x(118) & x(119) & x(131) & x(135) & x(138) & x(140) & x(141) & x(143) & x(151) & x(164) & x(187) & x(191) & x(193) & x(197) & x(213) & x(214) & x(221) & x(222) & x(235) & x(241) & x(243) & x(254);
    y(111) <= not(p111_out);
    p111 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00011110000001100100111100101001100011000",
            TABLE => "01111111000101110001011100000001000101110000000100000001000000000111111000010111000101111000000100010111100000011000000111101000011010011001011010010110011010011001011001101001011010011001011011101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011001000000110101001101010011111101000000000100000001000000110101000100001011010100110101001011110100101011010000100100001011010100011010011001011010010110011010011001011001101001011010011001011000010111011111110000000100010111000000010001011100000000000000010001011101111110100000010001011110000001000101111110100010000001100101100110100101101001100101100110100110010110100101100110100110110010111110110010000010110010001000001011001000000000001000001011001011011011001001001011001000100100101100100100110100100100100101100110100101101001100101100110100110010110100101100110100110000000111010001110100011111110000000001000000010000000111010001000000111101000111010000111111000010111100000011000000111101000100101100110100101101001100101100110100110010110100101100110100110000000111010001110100011111110100000011110100011101000011111101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p111_in,
            y(0) => p111_out,
            y(1 to 14 - 1) => dummy111
        );


    p112_in <= x(6) & x(10) & x(14) & x(16) & x(43) & x(53) & x(54) & x(66) & x(74) & x(76) & x(81) & x(99) & x(119) & x(128) & x(130) & x(140) & x(150) & x(156) & x(168) & x(182) & x(186) & x(207) & x(209) & x(214) & x(245) & x(250);
    y(112) <= not(p112_out);
    p112 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11110010111000110000111100",
            TABLE => "000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p112_in,
            y(0) => p112_out,
            y(1 to 14 - 1) => dummy112
        );


    p113_in <= x(5) & x(16) & x(25) & x(30) & x(48) & x(53) & x(56) & x(59) & x(62) & x(70) & x(76) & x(89) & x(92) & x(107) & x(110) & x(111) & x(113) & x(122) & x(124) & x(137) & x(142) & x(161) & x(166) & x(169) & x(179) & x(180) & x(182) & x(193) & x(197) & x(198) & x(211) & x(218) & x(229) & x(232) & x(236) & x(247) & x(252) & x(255);
    y(113) <= not(p113_out);
    p113 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110011011011010011011011010010011000",
            TABLE => "000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 4,
            B => -16,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p113_in,
            y(0) => p113_out,
            y(1 to 15 - 1) => dummy113
        );


    p114_in <= x(44) & x(47) & x(50) & x(60) & x(61) & x(68) & x(82) & x(86) & x(90) & x(95) & x(97) & x(98) & x(106) & x(111) & x(112) & x(113) & x(132) & x(134) & x(151) & x(154) & x(161) & x(162) & x(187) & x(191) & x(192) & x(195) & x(196) & x(203) & x(207) & x(221) & x(236) & x(239) & x(244) & x(247);
    y(114) <= not(p114_out);
    p114 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100110100011100101110100100111000",
            TABLE => "0111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101101101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010010010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101100000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010010111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101101000000011101000100000011110100010010110011010010000000000000000",
            SHIFT => 3,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p114_in,
            y(0) => p114_out,
            y(1 to 14 - 1) => dummy114
        );


    p115_in <= x(4) & x(27) & x(31) & x(36) & x(52) & x(66) & x(71) & x(77) & x(93) & x(96) & x(156) & x(167) & x(175) & x(176) & x(178) & x(179) & x(182) & x(192) & x(201) & x(220) & x(252);
    y(115) <= not(p115_out);
    p115 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100011001000000000111",
            TABLE => "011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 4,
            B => 7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p115_in,
            y(0) => p115_out,
            y(1 to 14 - 1) => dummy115
        );


    p116_in <= x(23) & x(32) & x(35) & x(49) & x(55) & x(58) & x(69) & x(73) & x(81) & x(109) & x(127) & x(156) & x(168) & x(171) & x(186) & x(195) & x(203) & x(204) & x(205) & x(241) & x(252);
    y(116) <= not(p116_out);
    p116 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011010011110011011100",
            TABLE => "001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001100011101001011011111111",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p116_in,
            y(0) => p116_out,
            y(1 to 14 - 1) => dummy116
        );


    p117_in <= x(3) & x(9) & x(13) & x(17) & x(26) & x(38) & x(52) & x(66) & x(68) & x(79) & x(87) & x(95) & x(110) & x(112) & x(126) & x(130) & x(135) & x(136) & x(140) & x(160) & x(162) & x(163) & x(176) & x(178) & x(179) & x(214) & x(218) & x(227) & x(230) & x(238) & x(243) & x(244) & x(253) & x(254);
    y(117) <= not(p117_out);
    p117 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001111110100001100000000001000010",
            TABLE => "0001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010011011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101101011001000100000101100100010010010010110011010010000000000000000",
            SHIFT => 3,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p117_in,
            y(0) => p117_out,
            y(1 to 14 - 1) => dummy117
        );


    p118_in <= x(4) & x(6) & x(9) & x(31) & x(66) & x(75) & x(83) & x(100) & x(123) & x(126) & x(130) & x(148) & x(151) & x(179) & x(199) & x(204) & x(211) & x(226) & x(232) & x(243) & x(250);
    y(118) <= not(p118_out);
    p118 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010101110101011010110",
            TABLE => "010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110001010110110100111111111",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p118_in,
            y(0) => p118_out,
            y(1 to 14 - 1) => dummy118
        );


    p119_in <= x(16) & x(18) & x(19) & x(26) & x(27) & x(40) & x(48) & x(77) & x(87) & x(102) & x(130) & x(147) & x(153) & x(154) & x(163) & x(179) & x(182) & x(183) & x(188) & x(200) & x(203) & x(213) & x(226) & x(228) & x(229) & x(234) & x(241) & x(243);
    y(119) <= not(p119_out);
    p119 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111000110100100000110110100",
            TABLE => "0000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101101110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101100001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010011000111000001000100011100001100010010110011010010000000000000000",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p119_in,
            y(0) => p119_out,
            y(1 to 14 - 1) => dummy119
        );


    p120_in <= x(4) & x(11) & x(20) & x(56) & x(87) & x(93) & x(122) & x(130) & x(143) & x(144) & x(147) & x(148) & x(153) & x(228) & x(243) & x(247);
    y(120) <= not(p120_out);
    p120 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110011000111011",
            TABLE => "0100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101100001000001110001000110000111000110010110011010010000000000000000",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p120_in,
            y(0) => p120_out,
            y(1 to 14 - 1) => dummy120
        );


    p121_in <= x(0) & x(2) & x(12) & x(20) & x(30) & x(38) & x(47) & x(48) & x(58) & x(60) & x(62) & x(64) & x(70) & x(81) & x(106) & x(108) & x(109) & x(116) & x(127) & x(132) & x(146) & x(156) & x(157) & x(170) & x(173) & x(187) & x(197) & x(198) & x(205) & x(219) & x(236) & x(238) & x(240) & x(241) & x(247);
    y(121) <= not(p121_out);
    p121 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101000100110010000010111000110010",
            TABLE => "10110010111110110010000010110010001000001011001000000000001000001011001011011011001001001011001000100100101100100100110100100100100101100110100101101001100101100110100110010110100101100110100111010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100110001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100111011111010011010100110100000100010011010000010000000100000000001101101101001101010011010010010001001101001001000010010010110010100101100110100101101001100101100110100110010110100101100110100101000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011010110010001000001111101110110010101100100010010011011011101100101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p121_in,
            y(0) => p121_out,
            y(1 to 14 - 1) => dummy121
        );


    p122_in <= x(4) & x(10) & x(26) & x(38) & x(54) & x(75) & x(84) & x(86) & x(107) & x(142) & x(162) & x(164) & x(174) & x(179) & x(182) & x(224) & x(233) & x(240) & x(248) & x(252);
    y(122) <= not(p122_out);
    p122 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01011101100001001110",
            TABLE => "000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 4,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p122_in,
            y(0) => p122_out,
            y(1 to 14 - 1) => dummy122
        );


    p123_in <= x(33) & x(51) & x(58) & x(64) & x(79) & x(81) & x(90) & x(103) & x(105) & x(106) & x(112) & x(128) & x(131) & x(132) & x(134) & x(140) & x(142) & x(153) & x(154) & x(166) & x(181) & x(186) & x(198) & x(213) & x(215) & x(218) & x(227) & x(231) & x(246);
    y(123) <= not(p123_out);
    p123 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11000101110001000111001100100",
            TABLE => "01000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011000001000100011101000111011101111000000000000100000001000100011100001100010001110100011101110011101110001000110000001100010001110011010011001011010010110011010011001011001101001011010011001011011010100010000001111110111010100010000000000000011010100010000001101010001000010101111011101010001000010001010111101010001000010100101100110100101101001100101100110100110010110100101100110100100010000000000000111000100010000011100010001000011110111011100010001100010001110011100010001100001110001000110001110011101110001100101100110100101101001100101100110100110010110100101100110100111101111100011101000111000001000111001111000111010001110000110000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 3,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p123_in,
            y(0) => p123_out,
            y(1 to 13 - 1) => dummy123
        );


    p124_in <= x(23) & x(26) & x(65) & x(69) & x(76) & x(78) & x(89) & x(91) & x(107) & x(116) & x(129) & x(157) & x(163) & x(182) & x(190) & x(192) & x(197) & x(211) & x(220) & x(226) & x(232) & x(234) & x(251) & x(252);
    y(124) <= not(p124_out);
    p124 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000010011011110101001000",
            TABLE => "111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p124_in,
            y(0) => p124_out,
            y(1 to 14 - 1) => dummy124
        );


    p125_in <= x(9) & x(19) & x(23) & x(39) & x(40) & x(43) & x(52) & x(82) & x(92) & x(97) & x(100) & x(129) & x(131) & x(145) & x(165) & x(191) & x(192) & x(211) & x(213) & x(225) & x(254);
    y(125) <= not(p125_out);
    p125 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011011100010110000001",
            TABLE => "000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001110101001001011011111111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p125_in,
            y(0) => p125_out,
            y(1 to 14 - 1) => dummy125
        );


    p126_in <= x(7) & x(18) & x(25) & x(30) & x(37) & x(39) & x(56) & x(59) & x(62) & x(75) & x(79) & x(87) & x(103) & x(118) & x(124) & x(163) & x(180) & x(207) & x(210) & x(218) & x(220) & x(235) & x(238) & x(242) & x(243) & x(246) & x(253);
    y(126) <= not(p126_out);
    p126 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100010001010100100110010110",
            TABLE => "101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110001010110110100111111111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p126_in,
            y(0) => p126_out,
            y(1 to 14 - 1) => dummy126
        );


    p127_in <= x(4) & x(19) & x(20) & x(27) & x(49) & x(54) & x(62) & x(63) & x(114) & x(139) & x(143) & x(147) & x(153) & x(179) & x(196) & x(239) & x(251);
    y(127) <= not(p127_out);
    p127 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00100100000111000",
            TABLE => "11010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100111111101110101001101010001000000110101000100000001000000000000001011110111010100110101000100001011010100010000100100001000101011011010011001011010010110011010011001011001101001011010011001011010000000111010001110100011111110100000011110100011101000011111101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p127_in,
            y(0) => p127_out,
            y(1 to 14 - 1) => dummy127
        );


    p128_in <= x(7) & x(18) & x(20) & x(30) & x(36) & x(39) & x(44) & x(48) & x(49) & x(59) & x(67) & x(78) & x(94) & x(105) & x(110) & x(134) & x(147) & x(148) & x(162) & x(168) & x(169) & x(179) & x(180) & x(193) & x(199) & x(209) & x(210) & x(215) & x(219) & x(224) & x(234) & x(235) & x(253);
    y(128) <= not(p128_out);
    p128 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010101001111100100010011100110111",
            TABLE => "010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => 3,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p128_in,
            y(0) => p128_out,
            y(1 to 14 - 1) => dummy128
        );


    p129_in <= x(0) & x(9) & x(25) & x(40) & x(42) & x(43) & x(91) & x(99) & x(115) & x(140) & x(145) & x(147) & x(164) & x(193) & x(200) & x(211) & x(247) & x(254);
    y(129) <= not(p129_out);
    p129 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100101010111000011",
            TABLE => "010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p129_in,
            y(0) => p129_out,
            y(1 to 14 - 1) => dummy129
        );


    p130_in <= x(58) & x(82) & x(98) & x(101) & x(102) & x(103) & x(113) & x(139) & x(175) & x(176) & x(188) & x(192) & x(228) & x(232) & x(252);
    y(130) <= not(p130_out);
    p130 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010101111101110",
            TABLE => "010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110001010110110100111111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p130_in,
            y(0) => p130_out,
            y(1 to 14 - 1) => dummy130
        );


    p131_in <= x(3) & x(15) & x(16) & x(26) & x(44) & x(45) & x(47) & x(73) & x(80) & x(114) & x(128) & x(135) & x(152) & x(158) & x(164) & x(168) & x(170) & x(200) & x(203) & x(212) & x(219) & x(222) & x(224) & x(227) & x(230) & x(240);
    y(131) <= not(p131_out);
    p131 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11110000111101111100110010",
            TABLE => "000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p131_in,
            y(0) => p131_out,
            y(1 to 14 - 1) => dummy131
        );


    p132_in <= x(4) & x(6) & x(10) & x(17) & x(24) & x(26) & x(30) & x(44) & x(66) & x(67) & x(78) & x(81) & x(88) & x(92) & x(93) & x(95) & x(96) & x(110) & x(129) & x(136) & x(145) & x(147) & x(159) & x(160) & x(163) & x(166) & x(174) & x(180) & x(181) & x(183) & x(189) & x(194) & x(209) & x(214) & x(217) & x(222) & x(229) & x(230) & x(235) & x(243) & x(250) & x(254);
    y(132) <= not(p132_out);
    p132 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011010010001000111111111110010011100110101",
            TABLE => "001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p132_in,
            y(0) => p132_out,
            y(1 to 14 - 1) => dummy132
        );


    p133_in <= x(6) & x(7) & x(26) & x(29) & x(31) & x(67) & x(80) & x(86) & x(99) & x(101) & x(117) & x(123) & x(133) & x(149) & x(162) & x(188) & x(194) & x(218) & x(230) & x(236);
    y(133) <= not(p133_out);
    p133 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11000001001101010101",
            TABLE => "100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p133_in,
            y(0) => p133_out,
            y(1 to 14 - 1) => dummy133
        );


    p134_in <= x(31) & x(47) & x(55) & x(68) & x(80) & x(84) & x(86) & x(98) & x(99) & x(117) & x(122) & x(123) & x(128) & x(130) & x(161) & x(177) & x(186) & x(189) & x(205) & x(227) & x(245);
    y(134) <= not(p134_out);
    p134 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100011001010100100001",
            TABLE => "011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001110101001001011011111111",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p134_in,
            y(0) => p134_out,
            y(1 to 14 - 1) => dummy134
        );


    p135_in <= x(4) & x(10) & x(16) & x(18) & x(46) & x(51) & x(75) & x(94) & x(102) & x(108) & x(119) & x(132) & x(144) & x(158) & x(162) & x(166) & x(173) & x(178) & x(182) & x(191) & x(207) & x(209) & x(234);
    y(135) <= not(p135_out);
    p135 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110011001011010000111",
            TABLE => "00001000100011101000111011101111000000000000100000001000100011100001100010001110100011101110011101110001000110000001100010001110011010011001011010010110011010011001011001101001011010011001011000100000000000001011001000100000101100100010000011111011101100100010010001001101101100100010010010110010001001001101101110110010011010011001011010010110011010011001011001101001011010011001011000001000000000001000111000001000100011100000100011101111100011100001100001110001100011100001100010001110000110001110011110001110011010011001011010010110011010011001011001101001011010011001011001111111000101110001011100000001011111100001011100010111100000010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p135_in,
            y(0) => p135_out,
            y(1 to 14 - 1) => dummy135
        );


    p136_in <= x(6) & x(10) & x(20) & x(39) & x(40) & x(54) & x(66) & x(76) & x(77) & x(80) & x(86) & x(91) & x(96) & x(127) & x(136) & x(156) & x(162) & x(168) & x(171) & x(178) & x(182) & x(183) & x(188) & x(210) & x(230) & x(236) & x(242) & x(249);
    y(136) <= not(p136_out);
    p136 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110110100101100001001110101",
            TABLE => "0000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101101011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010011000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010100110100000100010011010010010001101001100101100000000000000000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p136_in,
            y(0) => p136_out,
            y(1 to 14 - 1) => dummy136
        );


    p137_in <= x(24) & x(26) & x(34) & x(55) & x(78) & x(86) & x(100) & x(103) & x(109) & x(117) & x(122) & x(155) & x(165) & x(196) & x(197) & x(198) & x(199) & x(201) & x(208) & x(212) & x(236) & x(252) & x(253);
    y(137) <= not(p137_out);
    p137 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01001000101010111110011",
            TABLE => "10110010001000001111101110110010001000000000000010110010001000001011001000100100110110111011001000100100010011011011001000100100100101100110100101101001100101100110100110010110100101100110100110110010111110110010000010110010001000001011001000000000001000001011001011011011001001001011001000100100101100100100110100100100100101100110100101101001100101100110100110010110100101100110100100000001000101110000000000000001000101110111111100000001000101111000000100010111111010001000000100010111011111101000000100010111011010011001011010010110011010011001011001101001011010011001011001110001000100001111011101110001011100010001100011100111011100010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p137_in,
            y(0) => p137_out,
            y(1 to 14 - 1) => dummy137
        );


    p138_in <= x(7) & x(16) & x(20) & x(41) & x(42) & x(48) & x(51) & x(58) & x(59) & x(60) & x(61) & x(64) & x(67) & x(70) & x(79) & x(80) & x(84) & x(89) & x(105) & x(113) & x(115) & x(123) & x(127) & x(133) & x(140) & x(144) & x(149) & x(160) & x(165) & x(166) & x(187) & x(192) & x(195) & x(197) & x(198) & x(201) & x(215) & x(217) & x(235) & x(241) & x(246) & x(254);
    y(138) <= not(p138_out);
    p138 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010100010001011001000100111100101000100111",
            TABLE => "100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p138_in,
            y(0) => p138_out,
            y(1 to 14 - 1) => dummy138
        );


    p139_in <= x(14) & x(53) & x(69) & x(70) & x(80) & x(86) & x(91) & x(99) & x(110) & x(115) & x(117) & x(119) & x(123) & x(128) & x(134) & x(152) & x(168) & x(194) & x(216) & x(222) & x(232) & x(236);
    y(139) <= not(p139_out);
    p139 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110101111010111110110",
            TABLE => "0010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101100000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p139_in,
            y(0) => p139_out,
            y(1 to 14 - 1) => dummy139
        );


    p140_in <= x(1) & x(4) & x(11) & x(17) & x(32) & x(36) & x(59) & x(75) & x(81) & x(117) & x(124) & x(137) & x(141) & x(143) & x(160) & x(167) & x(176) & x(179) & x(188) & x(192) & x(194) & x(201) & x(230) & x(245) & x(247) & x(249);
    y(140) <= not(p140_out);
    p140 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10101111100000111111101110",
            TABLE => "000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p140_in,
            y(0) => p140_out,
            y(1 to 14 - 1) => dummy140
        );


    p141_in <= x(11) & x(17) & x(29) & x(36) & x(40) & x(42) & x(57) & x(67) & x(70) & x(80) & x(120) & x(127) & x(129) & x(156) & x(177) & x(178) & x(179) & x(220) & x(227) & x(230) & x(245);
    y(141) <= not(p141_out);
    p141 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010011110001000001100",
            TABLE => "011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110100011101001011011111111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p141_in,
            y(0) => p141_out,
            y(1 to 14 - 1) => dummy141
        );


    p142_in <= x(5) & x(12) & x(15) & x(16) & x(58) & x(70) & x(74) & x(83) & x(87) & x(88) & x(89) & x(93) & x(104) & x(107) & x(108) & x(111) & x(118) & x(136) & x(166) & x(170) & x(172) & x(183) & x(186) & x(202) & x(210) & x(215) & x(218) & x(233) & x(234) & x(240) & x(244) & x(245) & x(246) & x(248) & x(249);
    y(142) <= not(p142_out);
    p142 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000001100000001110100000000111010",
            TABLE => "11101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011010000000111010001110100011111110000000001000000010000000111010001000000111101000111010000111111000010111100000011000000111101000100101100110100101101001100101100110100110010110100101100110100111110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100110000000111010000000000010000000111010001111111010000000111010001000000111101000000101111000000111101000011111101000000111101000100101100110100101101001100101100110100110010110100101100110100111111101110101001101010001000000110101000100000001000000000000001011110111010100110101000100001011010100010000100100001000101011011010011001011010010110011010011001011001101001011010011001011000100000101100101011001011111011001001001011001010110010110110110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p142_in,
            y(0) => p142_out,
            y(1 to 15 - 1) => dummy142
        );


    p143_in <= x(0) & x(1) & x(6) & x(11) & x(25) & x(39) & x(40) & x(43) & x(49) & x(50) & x(66) & x(78) & x(90) & x(91) & x(92) & x(100) & x(105) & x(110) & x(112) & x(134) & x(137) & x(147) & x(148) & x(159) & x(169) & x(178) & x(180) & x(189) & x(193) & x(204) & x(255);
    y(143) <= not(p143_out);
    p143 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000110011111110001110000111110",
            TABLE => "1111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p143_in,
            y(0) => p143_out,
            y(1 to 14 - 1) => dummy143
        );


    p144_in <= x(1) & x(21) & x(26) & x(51) & x(52) & x(58) & x(60) & x(66) & x(71) & x(83) & x(85) & x(95) & x(103) & x(127) & x(131) & x(192) & x(198) & x(213) & x(216) & x(243) & x(250);
    y(144) <= not(p144_out);
    p144 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000100100101010111010",
            TABLE => "111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001101100101001011011111111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p144_in,
            y(0) => p144_out,
            y(1 to 14 - 1) => dummy144
        );


    p145_in <= x(22) & x(28) & x(56) & x(57) & x(60) & x(66) & x(76) & x(82) & x(83) & x(97) & x(100) & x(103) & x(108) & x(117) & x(123) & x(124) & x(130) & x(135) & x(142) & x(154) & x(162) & x(165) & x(172) & x(173) & x(192) & x(198) & x(213) & x(215) & x(216) & x(231) & x(237) & x(245);
    y(145) <= not(p145_out);
    p145 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10101011111000010101010011110010",
            TABLE => "001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 3,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p145_in,
            y(0) => p145_out,
            y(1 to 14 - 1) => dummy145
        );


    p146_in <= x(2) & x(8) & x(14) & x(22) & x(30) & x(42) & x(44) & x(50) & x(64) & x(67) & x(69) & x(75) & x(77) & x(81) & x(92) & x(105) & x(122) & x(139) & x(141) & x(145) & x(160) & x(162) & x(164) & x(170) & x(173) & x(177) & x(183) & x(193) & x(197) & x(211) & x(213) & x(219) & x(232) & x(239) & x(245) & x(247);
    y(146) <= not(p146_out);
    p146 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000111011110001001100011101101111100",
            TABLE => "011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p146_in,
            y(0) => p146_out,
            y(1 to 14 - 1) => dummy146
        );


    p147_in <= x(4) & x(47) & x(58) & x(60) & x(70) & x(73) & x(82) & x(83) & x(89) & x(95) & x(109) & x(113) & x(115) & x(117) & x(123) & x(126) & x(129) & x(131) & x(151) & x(163) & x(191) & x(192) & x(211) & x(216) & x(236) & x(239) & x(243) & x(250);
    y(147) <= not(p147_out);
    p147 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110110010000110011000011001",
            TABLE => "0000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101101110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101101101010001000000010000000000000011111101110101001101010001000000110101000100001001000010001010111011110111010100110101000100001010010110011010010110100110010110011010011001011010010110011010010100000011010100010000101101010001101001100101100000000000000000",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p147_in,
            y(0) => p147_out,
            y(1 to 13 - 1) => dummy147
        );


    p148_in <= x(19) & x(37) & x(38) & x(48) & x(59) & x(71) & x(84) & x(100) & x(101) & x(124) & x(130) & x(188) & x(208) & x(222) & x(228) & x(255);
    y(148) <= not(p148_out);
    p148 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010101101011010",
            TABLE => "0010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101100000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010010000010110010001001001011001001101001100101100000000000000000",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p148_in,
            y(0) => p148_out,
            y(1 to 14 - 1) => dummy148
        );


    p149_in <= x(4) & x(6) & x(8) & x(10) & x(21) & x(34) & x(44) & x(53) & x(63) & x(96) & x(97) & x(101) & x(102) & x(104) & x(110) & x(129) & x(133) & x(143) & x(144) & x(147) & x(153) & x(163) & x(164) & x(171) & x(172) & x(173) & x(174) & x(183) & x(184) & x(193) & x(199) & x(214) & x(233) & x(248);
    y(149) <= not(p149_out);
    p149 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000110000011100110000101111110000",
            TABLE => "0111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101101111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 3,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p149_in,
            y(0) => p149_out,
            y(1 to 14 - 1) => dummy149
        );


    p150_in <= x(4) & x(6) & x(7) & x(8) & x(17) & x(21) & x(26) & x(37) & x(39) & x(59) & x(62) & x(66) & x(75) & x(88) & x(96) & x(126) & x(130) & x(135) & x(143) & x(156) & x(169) & x(187) & x(191) & x(197) & x(200) & x(248) & x(249) & x(252) & x(255);
    y(150) <= not(p150_out);
    p150 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10001111101101001110100110011",
            TABLE => "01110001000100000001000000000000111101110111000101110001000100000111000100011000000110001000111011100111011100010111000100011000011010011001011010010110011010011001011001101001011010011001011000000000000100000001000001110001000100000111000101110001111101111000111000011000000110000111000100011000011100010111000111100111011010011001011010010110011010011001011001101001011010011001011001110001000100001111011101110001000100000000000001110001000100000111000100011000111001110111000100011000100011100111000100011000011010011001011010010110011010011001011001101001011010011001011001000000110101000000000001000000110101001111110101000000110101000100001011010100001010110100001011010100101111010100001011010100011010011001011010010110011010011001011001101001011010011001011001110001000100001111011101110001011100010001100011100111011100010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p150_in,
            y(0) => p150_out,
            y(1 to 14 - 1) => dummy150
        );


    p151_in <= x(3) & x(18) & x(20) & x(42) & x(54) & x(62) & x(66) & x(74) & x(76) & x(82) & x(83) & x(101) & x(103) & x(106) & x(128) & x(141) & x(160) & x(189) & x(196) & x(197) & x(207) & x(216) & x(219) & x(234) & x(249) & x(251);
    y(151) <= not(p151_out);
    p151 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000110000110100011011001",
            TABLE => "110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p151_in,
            y(0) => p151_out,
            y(1 to 14 - 1) => dummy151
        );


    p152_in <= x(2) & x(5) & x(7) & x(26) & x(32) & x(34) & x(54) & x(64) & x(65) & x(69) & x(81) & x(102) & x(108) & x(126) & x(137) & x(152) & x(156) & x(166) & x(168) & x(171) & x(173) & x(178) & x(184) & x(197) & x(200) & x(205) & x(208) & x(245);
    y(152) <= not(p152_out);
    p152 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000010111011111101011100010",
            TABLE => "1111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010011011001000100000101100100010010010010110011010010000000000000000",
            SHIFT => 3,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p152_in,
            y(0) => p152_out,
            y(1 to 13 - 1) => dummy152
        );


    p153_in <= x(1) & x(14) & x(17) & x(18) & x(19) & x(21) & x(33) & x(35) & x(36) & x(60) & x(72) & x(78) & x(89) & x(123) & x(132) & x(149) & x(167) & x(182) & x(192) & x(213) & x(217) & x(232) & x(248);
    y(153) <= not(p153_out);
    p153 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11011100101111011100100",
            TABLE => "00000001000000000001011100000001000101110000000101111111000101111000000111101000000101111000000100010111100000010111111000010111011010011001011010010110011010011001011001101001011010011001011001110001111101110001000001110001000100000111000100000000000100000111000111100111000110000111000100011000011100011000111000011000011010011001011010010110011010011001011001101001011010011001011000000001000000000001011100000001000101110000000101111111000101111000000111101000000101111000000100010111100000010111111000010111011010011001011010010110011010011001011001101001011010011001011011101111100011101000111000001000111001111000111010001110000110000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p153_in,
            y(0) => p153_out,
            y(1 to 14 - 1) => dummy153
        );


    p154_in <= x(8) & x(14) & x(21) & x(27) & x(44) & x(63) & x(105) & x(106) & x(127) & x(135) & x(136) & x(144) & x(161) & x(164) & x(182) & x(185) & x(203) & x(210) & x(211) & x(212) & x(215) & x(223) & x(225) & x(232) & x(242) & x(255);
    y(154) <= not(p154_out);
    p154 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00110011110011100110001101",
            TABLE => "100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p154_in,
            y(0) => p154_out,
            y(1 to 14 - 1) => dummy154
        );


    p155_in <= x(12) & x(39) & x(47) & x(50) & x(51) & x(68) & x(80) & x(82) & x(90) & x(98) & x(114) & x(115) & x(118) & x(126) & x(128) & x(132) & x(151) & x(158) & x(187) & x(188) & x(221) & x(227);
    y(155) <= not(p155_out);
    p155 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010110001001001101111",
            TABLE => "0001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010011110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p155_in,
            y(0) => p155_out,
            y(1 to 14 - 1) => dummy155
        );


    p156_in <= x(8) & x(27) & x(62) & x(82) & x(98) & x(104) & x(139) & x(153) & x(176) & x(187) & x(203) & x(205) & x(216) & x(218) & x(236) & x(244) & x(255);
    y(156) <= not(p156_out);
    p156 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10001001011010100",
            TABLE => "10110010001000000010000000000000111110111011001010110010001000001011001000100100001001000100110111011011101100101011001000100100100101100110100101101001100101100110100110010110100101100110100100101011000000101011111100101011000000100000000000101011000000100010101101000010101111010010101101000010110101000010101101000010011010011001011010010110011010011001011001101001011010011001011010001110000010001110111110001110100011100001100011100111100011101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p156_in,
            y(0) => p156_out,
            y(1 to 14 - 1) => dummy156
        );


    p157_in <= x(2) & x(13) & x(34) & x(37) & x(45) & x(61) & x(69) & x(83) & x(90) & x(103) & x(114) & x(126) & x(133) & x(137) & x(152) & x(171) & x(178) & x(194) & x(195) & x(196) & x(200) & x(223) & x(225) & x(233) & x(249) & x(255);
    y(157) <= not(p157_out);
    p157 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10010100011000010001101101",
            TABLE => "010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 3,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p157_in,
            y(0) => p157_out,
            y(1 to 13 - 1) => dummy157
        );


    p158_in <= x(8) & x(12) & x(20) & x(61) & x(62) & x(64) & x(67) & x(74) & x(79) & x(81) & x(83) & x(86) & x(94) & x(103) & x(105) & x(106) & x(127) & x(128) & x(135) & x(140) & x(145) & x(157) & x(160) & x(161) & x(164) & x(183) & x(185) & x(200) & x(214) & x(223) & x(242) & x(254);
    y(158) <= not(p158_out);
    p158 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11000100101010000101101000101111",
            TABLE => "010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 3,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p158_in,
            y(0) => p158_out,
            y(1 to 14 - 1) => dummy158
        );


    p159_in <= x(1) & x(11) & x(43) & x(52) & x(56) & x(71) & x(75) & x(79) & x(85) & x(89) & x(91) & x(92) & x(98) & x(99) & x(116) & x(119) & x(132) & x(141) & x(145) & x(151) & x(159) & x(168) & x(170) & x(177) & x(185) & x(186) & x(189) & x(200) & x(209) & x(219) & x(223) & x(225) & x(237);
    y(159) <= not(p159_out);
    p159 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000010101101011011010011110011",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001011100010110100111111111",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p159_in,
            y(0) => p159_out,
            y(1 to 15 - 1) => dummy159
        );


    p160_in <= x(14) & x(28) & x(62) & x(148) & x(158) & x(166) & x(238) & x(247);
    y(160) <= not(p160_out);
    p160 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11100011",
            TABLE => "000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 5,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p160_in,
            y(0) => p160_out,
            y(1 to 14 - 1) => dummy160
        );


    p161_in <= x(0) & x(1) & x(4) & x(6) & x(8) & x(21) & x(44) & x(45) & x(48) & x(53) & x(70) & x(83) & x(88) & x(92) & x(109) & x(110) & x(121) & x(122) & x(138) & x(152) & x(156) & x(164) & x(173) & x(186) & x(194) & x(204) & x(216) & x(226) & x(236) & x(250) & x(252);
    y(161) <= not(p161_out);
    p161 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010010000101100001011110111110",
            TABLE => "1101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101101000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p161_in,
            y(0) => p161_out,
            y(1 to 15 - 1) => dummy161
        );


    p162_in <= x(22) & x(32) & x(37) & x(39) & x(44) & x(49) & x(63) & x(65) & x(67) & x(77) & x(83) & x(125) & x(131) & x(133) & x(143) & x(173) & x(179) & x(183) & x(196) & x(201) & x(244);
    y(162) <= not(p162_out);
    p162 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011111100100101000100",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001100011101001011011111111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p162_in,
            y(0) => p162_out,
            y(1 to 14 - 1) => dummy162
        );


    p163_in <= x(15) & x(21) & x(26) & x(28) & x(40) & x(47) & x(57) & x(62) & x(88) & x(96) & x(104) & x(112) & x(118) & x(121) & x(151) & x(162) & x(164) & x(172) & x(175) & x(176) & x(187) & x(209) & x(231) & x(248) & x(253);
    y(163) <= not(p163_out);
    p163 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111001110110001111101100",
            TABLE => "0000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p163_in,
            y(0) => p163_out,
            y(1 to 13 - 1) => dummy163
        );


    p164_in <= x(10) & x(12) & x(14) & x(16) & x(18) & x(21) & x(36) & x(51) & x(66) & x(74) & x(78) & x(86) & x(99) & x(101) & x(114) & x(152) & x(161) & x(162) & x(174) & x(199) & x(201) & x(202) & x(205) & x(209) & x(233) & x(251);
    y(164) <= not(p164_out);
    p164 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10011110010100101000011111",
            TABLE => "000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p164_in,
            y(0) => p164_out,
            y(1 to 14 - 1) => dummy164
        );


    p165_in <= x(3) & x(4) & x(6) & x(8) & x(30) & x(63) & x(84) & x(93) & x(95) & x(96) & x(102) & x(104) & x(121) & x(122) & x(129) & x(133) & x(146) & x(155) & x(163) & x(169) & x(196) & x(208) & x(224) & x(226) & x(233) & x(235) & x(244);
    y(165) <= not(p165_out);
    p165 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101111000100101000101000100",
            TABLE => "000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001100011101001011011111111",
            SHIFT => 3,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p165_in,
            y(0) => p165_out,
            y(1 to 13 - 1) => dummy165
        );


    p166_in <= x(4) & x(7) & x(10) & x(14) & x(40) & x(50) & x(52) & x(68) & x(86) & x(88) & x(90) & x(101) & x(112) & x(130) & x(134) & x(162) & x(176) & x(177) & x(178) & x(191) & x(195) & x(203) & x(222) & x(232) & x(250) & x(254);
    y(166) <= not(p166_out);
    p166 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10010100011111111111011110",
            TABLE => "010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 4,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p166_in,
            y(0) => p166_out,
            y(1 to 14 - 1) => dummy166
        );


    p167_in <= x(27) & x(65) & x(93) & x(97) & x(117) & x(132) & x(142) & x(160) & x(169) & x(230) & x(236);
    y(167) <= not(p167_out);
    p167 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10010011010",
            TABLE => "10001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100100100000101100101011001011111011001001001011001010110010110110110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p167_in,
            y(0) => p167_out,
            y(1 to 14 - 1) => dummy167
        );


    p168_in <= x(3) & x(13) & x(14) & x(25) & x(30) & x(38) & x(39) & x(45) & x(59) & x(107) & x(140) & x(156) & x(165) & x(169) & x(201) & x(210) & x(214) & x(215) & x(216) & x(228) & x(229) & x(238) & x(251);
    y(168) <= not(p168_out);
    p168 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10011110110100000111001",
            TABLE => "00010111000000010000000100000000011111110001011100010111000000010001011110000001100000011110100001111110000101110001011110000001100101100110100101101001100101100110100110010110100101100110100100000100010011010000000000000100010011011101111100000100010011010010010001001101101100100010010001001101110110110010010001001101100101100110100101101001100101100110100110010110100101100110100111111101110101001101010001000000110101000100000001000000000000001011110111010100110101000100001011010100010000100100001000101011011010011001011010010110011010011001011001101001011010011001011001000000110101001101010011111101010000101101010011010100101111010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -14,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p168_in,
            y(0) => p168_out,
            y(1 to 14 - 1) => dummy168
        );


    p169_in <= x(11) & x(14) & x(19) & x(37) & x(53) & x(60) & x(75) & x(83) & x(85) & x(95) & x(121) & x(129) & x(133) & x(158) & x(196) & x(205) & x(212) & x(215) & x(216) & x(225) & x(226) & x(231) & x(242);
    y(169) <= not(p169_out);
    p169 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00011000101101101011000",
            TABLE => "10111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100101110001111101110001000001110001000100000111000100000000000100000111000111100111000110000111000100011000011100011000111000011000011010011001011010010110011010011001011001101001011010011001011000100000101100101011001011111011000000000010000000100000101100100010010010110010101100101101101101001101001001000010010010110010011010011001011010010110011010011001011001101001011010011001011010000000111010001110100011111110100000011110100011101000011111101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p169_in,
            y(0) => p169_out,
            y(1 to 14 - 1) => dummy169
        );


    p170_in <= x(4) & x(20) & x(34) & x(49) & x(56) & x(58) & x(74) & x(88) & x(89) & x(100) & x(101) & x(103) & x(106) & x(107) & x(126) & x(161) & x(165) & x(179) & x(181) & x(213) & x(218) & x(250) & x(254);
    y(170) <= not(p170_out);
    p170 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10010100100000001010111",
            TABLE => "01001101000001000000010000000000110111110100110101001101000001000100110100100100001001001011001011011011010011010100110100100100011010011001011010010110011010011001011001101001011010011001011011101000111111101000000011101000100000001110100000000000100000001110100001111110100000011110100010000001111010000001011110000001011010011001011010010110011010011001011001101001011010011001011011111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011000010111000000010111111100010111000101111000000101111110000101111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p170_in,
            y(0) => p170_out,
            y(1 to 14 - 1) => dummy170
        );


    p171_in <= x(4) & x(23) & x(31) & x(35) & x(47) & x(55) & x(73) & x(80) & x(83) & x(89) & x(117) & x(126) & x(128) & x(166) & x(168) & x(171) & x(172) & x(186) & x(194) & x(199) & x(204) & x(225) & x(234) & x(243) & x(255);
    y(171) <= not(p171_out);
    p171 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110000110011110001100110",
            TABLE => "1000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p171_in,
            y(0) => p171_out,
            y(1 to 14 - 1) => dummy171
        );


    p172_in <= x(9) & x(39) & x(50) & x(59) & x(78) & x(82) & x(85) & x(100) & x(105) & x(109) & x(112) & x(113) & x(130) & x(132) & x(134) & x(151) & x(187) & x(195) & x(203) & x(204) & x(210) & x(216) & x(222) & x(243);
    y(172) <= not(p172_out);
    p172 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000100111000010111000100",
            TABLE => "111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p172_in,
            y(0) => p172_out,
            y(1 to 13 - 1) => dummy172
        );


    p173_in <= x(11) & x(17) & x(23) & x(29) & x(30) & x(37) & x(39) & x(45) & x(50) & x(52) & x(63) & x(95) & x(101) & x(130) & x(133) & x(139) & x(140) & x(141) & x(160) & x(188) & x(207) & x(217) & x(225) & x(249);
    y(173) <= not(p173_out);
    p173 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101100010101001010111100",
            TABLE => "000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p173_in,
            y(0) => p173_out,
            y(1 to 13 - 1) => dummy173
        );


    p174_in <= x(8) & x(26) & x(29) & x(34) & x(37) & x(41) & x(46) & x(47) & x(59) & x(62) & x(76) & x(80) & x(82) & x(83) & x(90) & x(91) & x(95) & x(98) & x(123) & x(126) & x(128) & x(130) & x(131) & x(171) & x(175) & x(194) & x(210) & x(216) & x(219) & x(224) & x(234) & x(243);
    y(174) <= not(p174_out);
    p174 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11001111010000000110011100110100",
            TABLE => "000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p174_in,
            y(0) => p174_out,
            y(1 to 15 - 1) => dummy174
        );


    p175_in <= x(11) & x(15) & x(29) & x(30) & x(31) & x(40) & x(41) & x(47) & x(80) & x(91) & x(98) & x(117) & x(127) & x(132) & x(145) & x(147) & x(162) & x(175) & x(183) & x(196) & x(221) & x(227) & x(236) & x(244) & x(247);
    y(175) <= not(p175_out);
    p175 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100011100111101001011100",
            TABLE => "1101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010010001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010010000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p175_in,
            y(0) => p175_out,
            y(1 to 14 - 1) => dummy175
        );


    p176_in <= x(4) & x(10) & x(16) & x(21) & x(24) & x(51) & x(54) & x(56) & x(57) & x(74) & x(75) & x(76) & x(96) & x(106) & x(108) & x(140) & x(144) & x(154) & x(160) & x(166) & x(167) & x(182) & x(198) & x(201) & x(209) & x(216) & x(224);
    y(176) <= not(p176_out);
    p176 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100001001000001000000101011",
            TABLE => "110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001011100010110100111111111",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p176_in,
            y(0) => p176_out,
            y(1 to 14 - 1) => dummy176
        );


    p177_in <= x(7) & x(30) & x(33) & x(37) & x(39) & x(49) & x(57) & x(77) & x(78) & x(87) & x(93) & x(100) & x(101) & x(103) & x(105) & x(130) & x(136) & x(154) & x(160) & x(182) & x(205) & x(212) & x(224);
    y(177) <= not(p177_out);
    p177 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000010001101100001111",
            TABLE => "11101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011001110001000100000001000000000000111101110111000101110001000100000111000100011000000110001000111011100111011100010111000100011000011010011001011010010110011010011001011001101001011010011001011010000000111010001110100011111110000000001000000010000000111010001000000111101000111010000111111000010111100000011000000111101000100101100110100101101001100101100110100110010110100101100110100100010111011111110000000100010111000101110111111010000001000101111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p177_in,
            y(0) => p177_out,
            y(1 to 14 - 1) => dummy177
        );


    p178_in <= x(6) & x(12) & x(15) & x(27) & x(39) & x(60) & x(70) & x(78) & x(83) & x(89) & x(90) & x(103) & x(108) & x(111) & x(116) & x(117) & x(136) & x(145) & x(153) & x(157) & x(182) & x(184) & x(187) & x(194) & x(197) & x(210) & x(220) & x(223) & x(225) & x(234) & x(251);
    y(178) <= not(p178_out);
    p178 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000110110100010110000011011011",
            TABLE => "1111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101100111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101101111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p178_in,
            y(0) => p178_out,
            y(1 to 15 - 1) => dummy178
        );


    p179_in <= x(7) & x(8) & x(12) & x(16) & x(17) & x(21) & x(26) & x(39) & x(40) & x(47) & x(55) & x(88) & x(89) & x(99) & x(104) & x(118) & x(121) & x(135) & x(143) & x(147) & x(151) & x(152) & x(158) & x(164) & x(172) & x(175) & x(182) & x(187) & x(190) & x(195) & x(200) & x(202) & x(204) & x(209) & x(227) & x(241) & x(255);
    y(179) <= not(p179_out);
    p179 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110000011000101100111000001110000110",
            TABLE => "0000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101101000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101100000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101101111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p179_in,
            y(0) => p179_out,
            y(1 to 14 - 1) => dummy179
        );


    p180_in <= x(4) & x(6) & x(10) & x(16) & x(17) & x(24) & x(37) & x(50) & x(56) & x(62) & x(65) & x(66) & x(67) & x(75) & x(76) & x(82) & x(96) & x(99) & x(100) & x(108) & x(109) & x(119) & x(160) & x(173) & x(182) & x(201) & x(206) & x(216) & x(224) & x(239) & x(248) & x(250);
    y(180) <= not(p180_out);
    p180 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000011011110000101010111111101",
            TABLE => "111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 3,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p180_in,
            y(0) => p180_out,
            y(1 to 14 - 1) => dummy180
        );


    p181_in <= x(4) & x(6) & x(8) & x(17) & x(18) & x(19) & x(20) & x(25) & x(26) & x(53) & x(65) & x(66) & x(83) & x(87) & x(110) & x(129) & x(133) & x(135) & x(143) & x(147) & x(153) & x(157) & x(163) & x(164) & x(174) & x(179) & x(180) & x(215) & x(217) & x(226) & x(230) & x(232) & x(235) & x(241) & x(251);
    y(181) <= not(p181_out);
    p181 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10011101101111001110000110111100101",
            TABLE => "00010111000000010000000100000000011111110001011100010111000000010001011110000001100000011110100001111110000101110001011110000001100101100110100101101001100101100110100110010110100101100110100100010000011100010111000111110111000000000001000000010000011100010001100001110001011100011110011110001110000110000001100001110001100101100110100101101001100101100110100110010110100101100110100100010000000000000111000100010000011100010001000011110111011100010001100010001110011100010001100001110001000110001110011101110001100101100110100101101001100101100110100110010110100101100110100111010100010000000100000000000000111111011101010011010100010000001101010001000010010000100010101110111101110101001101010001000010100101100110100101101001100101100110100110010110100101100110100100000001000101110000000000000001000101110111111100000001000101111000000100010111111010001000000100010111011111101000000100010111011010011001011010010110011010011001011001101001011010011001011011011111010011010100110100000100110110110100110101001101001001001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p181_in,
            y(0) => p181_out,
            y(1 to 14 - 1) => dummy181
        );


    p182_in <= x(0) & x(1) & x(7) & x(8) & x(25) & x(32) & x(39) & x(40) & x(50) & x(53) & x(63) & x(77) & x(82) & x(102) & x(112) & x(122) & x(134) & x(147) & x(153) & x(169) & x(186) & x(189) & x(193) & x(203) & x(204) & x(206) & x(211) & x(228) & x(230) & x(232) & x(254);
    y(182) <= not(p182_out);
    p182 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000111010111010100011111011010",
            TABLE => "1111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010010010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 3,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p182_in,
            y(0) => p182_out,
            y(1 to 14 - 1) => dummy182
        );


    p183_in <= x(4) & x(14) & x(16) & x(40) & x(47) & x(50) & x(55) & x(56) & x(62) & x(74) & x(75) & x(76) & x(87) & x(88) & x(100) & x(107) & x(111) & x(112) & x(119) & x(130) & x(137) & x(147) & x(153) & x(156) & x(158) & x(163) & x(165) & x(167) & x(171) & x(176) & x(179) & x(195) & x(196) & x(198) & x(205) & x(231) & x(234) & x(247) & x(255);
    y(183) <= not(p183_out);
    p183 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001100010111011110101111110100110000100",
            TABLE => "100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001100011101001011011111111",
            SHIFT => 3,
            B => -13,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p183_in,
            y(0) => p183_out,
            y(1 to 14 - 1) => dummy183
        );


    p184_in <= x(1) & x(5) & x(10) & x(14) & x(20) & x(25) & x(37) & x(59) & x(62) & x(66) & x(68) & x(86) & x(100) & x(101) & x(105) & x(122) & x(130) & x(166) & x(177) & x(188) & x(206) & x(215) & x(228) & x(245) & x(247) & x(251) & x(255);
    y(184) <= not(p184_out);
    p184 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110110101100010111101001101",
            TABLE => "000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110010011010110100111111111",
            SHIFT => 4,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p184_in,
            y(0) => p184_out,
            y(1 to 14 - 1) => dummy184
        );


    p185_in <= x(4) & x(6) & x(10) & x(47) & x(48) & x(65) & x(76) & x(80) & x(85) & x(102) & x(108) & x(110) & x(114) & x(133) & x(150) & x(158) & x(166) & x(173) & x(208) & x(224) & x(249);
    y(185) <= not(p185_out);
    p185 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100101000110011001111",
            TABLE => "010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p185_in,
            y(0) => p185_out,
            y(1 to 14 - 1) => dummy185
        );


    p186_in <= x(3) & x(5) & x(16) & x(20) & x(27) & x(28) & x(30) & x(78) & x(80) & x(85) & x(86) & x(104) & x(111) & x(127) & x(148) & x(150) & x(161) & x(172) & x(173) & x(183) & x(184) & x(188) & x(189) & x(196) & x(199) & x(209) & x(210) & x(232) & x(238) & x(248) & x(253);
    y(186) <= not(p186_out);
    p186 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100001111000001000000011000011",
            TABLE => "1000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010011110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101101111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101101101010001000000010000000000000011111101110101001101010001000000110101000100001001000010001010111011110111010100110101000100001010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p186_in,
            y(0) => p186_out,
            y(1 to 14 - 1) => dummy186
        );


    p187_in <= x(13) & x(39) & x(47) & x(50) & x(70) & x(105) & x(113) & x(116) & x(130) & x(134) & x(135) & x(136) & x(140) & x(151) & x(154) & x(187) & x(216) & x(222) & x(236) & x(239) & x(249);
    y(187) <= not(p187_out);
    p187 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001011000000111110101",
            TABLE => "011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110010011010110100111111111",
            SHIFT => 4,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p187_in,
            y(0) => p187_out,
            y(1 to 14 - 1) => dummy187
        );


    p188_in <= x(2) & x(5) & x(27) & x(54) & x(69) & x(80) & x(93) & x(104) & x(108) & x(111) & x(131) & x(134) & x(137) & x(141) & x(152) & x(161) & x(180) & x(189) & x(193) & x(196) & x(201) & x(208) & x(214) & x(245) & x(247) & x(249) & x(255);
    y(188) <= not(p188_out);
    p188 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001110011101111111101110010",
            TABLE => "001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001101100101001011011111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p188_in,
            y(0) => p188_out,
            y(1 to 14 - 1) => dummy188
        );


    p189_in <= x(10) & x(12) & x(17) & x(22) & x(28) & x(31) & x(46) & x(58) & x(62) & x(64) & x(68) & x(74) & x(77) & x(97) & x(99) & x(103) & x(113) & x(138) & x(143) & x(154) & x(156) & x(161) & x(164) & x(178) & x(179) & x(191) & x(197) & x(205) & x(224) & x(243) & x(244) & x(249) & x(254);
    y(189) <= not(p189_out);
    p189 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010111100100011010001001110011101",
            TABLE => "000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001010011010110100111111111",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p189_in,
            y(0) => p189_out,
            y(1 to 14 - 1) => dummy189
        );


    p190_in <= x(3) & x(7) & x(13) & x(20) & x(22) & x(36) & x(47) & x(48) & x(54) & x(80) & x(85) & x(89) & x(107) & x(114) & x(119) & x(127) & x(145) & x(153) & x(156) & x(158) & x(168) & x(169) & x(172) & x(183) & x(185) & x(188) & x(189) & x(196) & x(198) & x(210) & x(219) & x(227) & x(237) & x(253);
    y(190) <= not(p190_out);
    p190 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111101110010001010001110110110110",
            TABLE => "0000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010010000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010011101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 3,
            B => 9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p190_in,
            y(0) => p190_out,
            y(1 to 14 - 1) => dummy190
        );


    p191_in <= x(14) & x(20) & x(40) & x(67) & x(86) & x(89) & x(101) & x(118) & x(120) & x(124) & x(130) & x(133) & x(144) & x(149) & x(151) & x(152) & x(159) & x(166) & x(168) & x(176) & x(177) & x(178) & x(199) & x(204) & x(217) & x(234) & x(241) & x(254);
    y(191) <= not(p191_out);
    p191 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101001110110011000111011000",
            TABLE => "0000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101100000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101101000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010011000000011101000100000011110100010010110011010010000000000000000",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p191_in,
            y(0) => p191_out,
            y(1 to 14 - 1) => dummy191
        );


    p192_in <= x(17) & x(53) & x(54) & x(55) & x(63) & x(72) & x(80) & x(91) & x(99) & x(100) & x(109) & x(119) & x(137) & x(156) & x(168) & x(172) & x(182) & x(186) & x(206) & x(209) & x(230) & x(232) & x(235) & x(237) & x(240) & x(241);
    y(192) <= not(p192_out);
    p192 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01001111100101101010100001",
            TABLE => "011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p192_in,
            y(0) => p192_out,
            y(1 to 14 - 1) => dummy192
        );


    p193_in <= x(0) & x(15) & x(19) & x(25) & x(41) & x(59) & x(63) & x(100) & x(103) & x(119) & x(152) & x(169) & x(174) & x(175) & x(186) & x(198) & x(203) & x(227) & x(228) & x(229) & x(234) & x(240) & x(251) & x(254);
    y(193) <= not(p193_out);
    p193 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001101111100011010101110",
            TABLE => "010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p193_in,
            y(0) => p193_out,
            y(1 to 14 - 1) => dummy193
        );


    p194_in <= x(12) & x(16) & x(22) & x(25) & x(26) & x(27) & x(30) & x(31) & x(39) & x(40) & x(58) & x(83) & x(89) & x(99) & x(102) & x(103) & x(130) & x(145) & x(152) & x(158) & x(161) & x(170) & x(185) & x(186) & x(189) & x(195) & x(199) & x(204) & x(207) & x(209) & x(223) & x(229) & x(233) & x(245);
    y(194) <= not(p194_out);
    p194 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111101010101001100111011001110010",
            TABLE => "0000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010010010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101100010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010011011001000100000101100100010010010010110011010010000000000000000",
            SHIFT => 4,
            B => 10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p194_in,
            y(0) => p194_out,
            y(1 to 15 - 1) => dummy194
        );


    p195_in <= x(3) & x(8) & x(31) & x(34) & x(37) & x(45) & x(51) & x(59) & x(61) & x(69) & x(85) & x(90) & x(92) & x(95) & x(96) & x(98) & x(100) & x(111) & x(125) & x(126) & x(133) & x(147) & x(155) & x(156) & x(180) & x(184) & x(188) & x(193) & x(203) & x(206) & x(232) & x(233) & x(235) & x(240);
    y(195) <= not(p195_out);
    p195 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100100010100011000001000000010100",
            TABLE => "0010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101101011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010011000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010011110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101101111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101101000111000001000100011100001100010010110011010010000000000000000",
            SHIFT => 3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p195_in,
            y(0) => p195_out,
            y(1 to 14 - 1) => dummy195
        );


    p196_in <= x(21) & x(26) & x(37) & x(40) & x(46) & x(57) & x(59) & x(62) & x(66) & x(69) & x(73) & x(97) & x(118) & x(119) & x(129) & x(135) & x(140) & x(160) & x(164) & x(167) & x(169) & x(174) & x(176) & x(177) & x(180) & x(182) & x(183) & x(185) & x(197) & x(202) & x(203) & x(212) & x(222) & x(223) & x(239) & x(242) & x(244) & x(248) & x(252);
    y(196) <= not(p196_out);
    p196 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000010100011101011000011100100110101110",
            TABLE => "111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001001010110110100111111111",
            SHIFT => 3,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p196_in,
            y(0) => p196_out,
            y(1 to 14 - 1) => dummy196
        );


    p197_in <= x(14) & x(110) & x(115) & x(129) & x(133) & x(151) & x(154) & x(159) & x(163) & x(166) & x(182) & x(192) & x(197) & x(208) & x(209) & x(211) & x(217) & x(221) & x(226) & x(232) & x(239) & x(253);
    y(197) <= not(p197_out);
    p197 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111000111110011000110",
            TABLE => "0000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101101000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p197_in,
            y(0) => p197_out,
            y(1 to 14 - 1) => dummy197
        );


    p198_in <= x(10) & x(32) & x(34) & x(44) & x(55) & x(60) & x(65) & x(67) & x(70) & x(81) & x(102) & x(113) & x(156) & x(168) & x(171) & x(184) & x(205) & x(216);
    y(198) <= not(p198_out);
    p198 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001000111010110101",
            TABLE => "111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p198_in,
            y(0) => p198_out,
            y(1 to 14 - 1) => dummy198
        );


    p199_in <= x(12) & x(17) & x(26) & x(46) & x(47) & x(48) & x(70) & x(92) & x(95) & x(98) & x(104) & x(109) & x(111) & x(115) & x(117) & x(131) & x(139) & x(142) & x(175) & x(209) & x(216) & x(244) & x(252) & x(255);
    y(199) <= not(p199_out);
    p199 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100110110100101010001000",
            TABLE => "001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -19,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p199_in,
            y(0) => p199_out,
            y(1 to 14 - 1) => dummy199
        );


    p200_in <= x(37) & x(48) & x(52) & x(54) & x(61) & x(64) & x(69) & x(79) & x(82) & x(83) & x(90) & x(95) & x(104) & x(126) & x(132) & x(134) & x(136) & x(140) & x(146) & x(156) & x(160) & x(178) & x(179) & x(203) & x(205) & x(234) & x(242) & x(243);
    y(200) <= not(p200_out);
    p200 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110100000000010001000001000",
            TABLE => "0000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101101110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101000000011101000100000011110100010010110011010010000000000000000",
            SHIFT => 3,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p200_in,
            y(0) => p200_out,
            y(1 to 13 - 1) => dummy200
        );


    p201_in <= x(8) & x(25) & x(28) & x(51) & x(52) & x(58) & x(67) & x(75) & x(84) & x(87) & x(89) & x(108) & x(110) & x(124) & x(133) & x(135) & x(136) & x(142) & x(149) & x(163) & x(178) & x(180) & x(193) & x(198) & x(206) & x(214) & x(218) & x(238) & x(246) & x(253) & x(254);
    y(201) <= not(p201_out);
    p201 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010010000111000111110001111101",
            TABLE => "0100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101101111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 3,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p201_in,
            y(0) => p201_out,
            y(1 to 14 - 1) => dummy201
        );


    p202_in <= x(0) & x(3) & x(5) & x(14) & x(15) & x(19) & x(20) & x(21) & x(28) & x(51) & x(58) & x(70) & x(73) & x(88) & x(105) & x(113) & x(118) & x(125) & x(132) & x(136) & x(144) & x(152) & x(158) & x(170) & x(175) & x(176) & x(179) & x(191) & x(193) & x(200) & x(212) & x(217) & x(219) & x(234) & x(235) & x(240);
    y(202) <= not(p202_out);
    p202 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010010010011010001001011001011001100",
            TABLE => "101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p202_in,
            y(0) => p202_out,
            y(1 to 15 - 1) => dummy202
        );


    p203_in <= x(23) & x(24) & x(71) & x(81) & x(83) & x(89) & x(99) & x(101) & x(120) & x(126) & x(128) & x(131) & x(152) & x(168) & x(171) & x(186) & x(188) & x(189) & x(194) & x(199) & x(205) & x(251) & x(254);
    y(203) <= not(p203_out);
    p203 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10101011011011000011011",
            TABLE => "00100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011000000010000000000010101100000010001010110000001010111111001010110100001011010100001010110100001000101011010000101011110100101011100101100110100101101001100101100110100110010110100101100110100110000000000000001110100010000000111010001000000011111110111010001000000100010111111010001000000111101000100000010111111011101000100101100110100101101001100101100110100110010110100101100110100100010000011100010111000111110111000110000111000101110001111001111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p203_in,
            y(0) => p203_out,
            y(1 to 14 - 1) => dummy203
        );


    p204_in <= x(1) & x(12) & x(14) & x(37) & x(43) & x(52) & x(55) & x(60) & x(64) & x(76) & x(82) & x(86) & x(92) & x(93) & x(112) & x(115) & x(126) & x(134) & x(137) & x(167) & x(168) & x(178) & x(186) & x(232) & x(237);
    y(204) <= not(p204_out);
    p204 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001110000010100000110000",
            TABLE => "0001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101101110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101101000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p204_in,
            y(0) => p204_out,
            y(1 to 14 - 1) => dummy204
        );


    p205_in <= x(16) & x(20) & x(21) & x(30) & x(47) & x(60) & x(70) & x(73) & x(88) & x(94) & x(107) & x(124) & x(128) & x(148) & x(165) & x(170) & x(179) & x(188) & x(198) & x(202) & x(219) & x(223) & x(226) & x(227) & x(241) & x(242) & x(247) & x(254);
    y(205) <= not(p205_out);
    p205 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100110100010010011001110110",
            TABLE => "0111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101101101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010011101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 3,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p205_in,
            y(0) => p205_out,
            y(1 to 13 - 1) => dummy205
        );


    p206_in <= x(2) & x(3) & x(4) & x(6) & x(13) & x(14) & x(27) & x(56) & x(59) & x(63) & x(65) & x(66) & x(69) & x(76) & x(78) & x(80) & x(85) & x(96) & x(101) & x(102) & x(105) & x(108) & x(114) & x(129) & x(134) & x(152) & x(154) & x(158) & x(173) & x(174) & x(192) & x(201) & x(212) & x(224) & x(233);
    y(206) <= not(p206_out);
    p206 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101110001110100011010011001101010",
            TABLE => "01110001111101110001000001110001000100000111000100000000000100000111000111100111000110000111000100011000011100011000111000011000011010011001011010010110011010011001011001101001011010011001011001110001000100000001000000000000111101110111000101110001000100000111000100011000000110001000111011100111011100010111000100011000011010011001011010010110011010011001011001101001011010011001011010000000111010000000000010000000111010001111111010000000111010001000000111101000000101111000000111101000011111101000000111101000100101100110100101101001100101100110100110010110100101100110100100001000000000001000111000001000100011100000100011101111100011100001100001110001100011100001100010001110000110001110011110001110011010011001011010010110011010011001011001101001011010011001011000010000000000000111000100010000011100010001000011110111011100010001100010001110011100010001100001110001000110001110011101110001100101100110100101101001100101100110100110010110100101100110100110110010111110110010000010110010101100101101101100100100101100101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p206_in,
            y(0) => p206_out,
            y(1 to 14 - 1) => dummy206
        );


    p207_in <= x(3) & x(31) & x(35) & x(43) & x(47) & x(51) & x(53) & x(68) & x(72) & x(80) & x(99) & x(101) & x(117) & x(119) & x(123) & x(128) & x(154) & x(156) & x(162) & x(171) & x(177) & x(180) & x(186) & x(189) & x(194) & x(230) & x(233) & x(236);
    y(207) <= not(p207_out);
    p207 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101011011110101011010001100",
            TABLE => "0000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101101000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010000100010001110000110001000111001101001100101100000000000000000",
            SHIFT => 3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p207_in,
            y(0) => p207_out,
            y(1 to 13 - 1) => dummy207
        );


    p208_in <= x(6) & x(11) & x(26) & x(30) & x(35) & x(38) & x(49) & x(50) & x(60) & x(63) & x(64) & x(75) & x(81) & x(84) & x(94) & x(104) & x(109) & x(132) & x(133) & x(141) & x(146) & x(149) & x(155) & x(156) & x(163) & x(169) & x(174) & x(196) & x(198) & x(209) & x(223) & x(226) & x(237) & x(239) & x(242) & x(244);
    y(208) <= not(p208_out);
    p208 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100101110110001000010101100100000100",
            TABLE => "010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p208_in,
            y(0) => p208_out,
            y(1 to 14 - 1) => dummy208
        );


    p209_in <= x(4) & x(10) & x(21) & x(28) & x(30) & x(34) & x(38) & x(42) & x(49) & x(51) & x(62) & x(68) & x(87) & x(99) & x(100) & x(112) & x(114) & x(118) & x(119) & x(125) & x(133) & x(139) & x(143) & x(144) & x(156) & x(161) & x(162) & x(177) & x(178) & x(188) & x(191) & x(201) & x(205) & x(215) & x(217) & x(224) & x(233) & x(234) & x(236) & x(239) & x(245) & x(247) & x(251);
    y(209) <= not(p209_out);
    p209 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110101110111010101001110100000011001101001",
            TABLE => "0010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101100000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101100001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010011110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101101000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 3,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p209_in,
            y(0) => p209_out,
            y(1 to 14 - 1) => dummy209
        );


    p210_in <= x(2) & x(4) & x(9) & x(20) & x(22) & x(23) & x(38) & x(44) & x(48) & x(74) & x(100) & x(101) & x(102) & x(119) & x(125) & x(144) & x(145) & x(173) & x(174) & x(183) & x(191) & x(203) & x(212) & x(213) & x(223) & x(225) & x(234) & x(251) & x(255);
    y(210) <= not(p210_out);
    p210 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01111000100110100111100101001",
            TABLE => "00000010001010110010101110111111000000000000001000000010001010110100001000101011001010111011110111010100010000100100001000101011100101100110100101101001100101100110100110010110100101100110100111010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100101000000110101000000000001000000110101001111110101000000110101000100001011010100001010110100001011010100101111010100001011010100011010011001011010010110011010011001011001101001011010011001011000000000010000000100000011010100010000001101010011010100111111010010101101000010010000101101010001000010110101001101010010111101100101100110100101101001100101100110100110010110100101100110100111010100111111010100000011010100110101001011110101000010110101001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p210_in,
            y(0) => p210_out,
            y(1 to 14 - 1) => dummy210
        );


    p211_in <= x(11) & x(17) & x(22) & x(36) & x(40) & x(44) & x(80) & x(98) & x(101) & x(103) & x(105) & x(126) & x(129) & x(132) & x(150) & x(162) & x(175) & x(181) & x(192) & x(202) & x(208) & x(212) & x(227) & x(232);
    y(211) <= not(p211_out);
    p211 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011010010000011000001010",
            TABLE => "001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p211_in,
            y(0) => p211_out,
            y(1 to 14 - 1) => dummy211
        );


    p212_in <= x(0) & x(3) & x(15) & x(20) & x(25) & x(30) & x(37) & x(48) & x(53) & x(59) & x(61) & x(62) & x(71) & x(77) & x(78) & x(90) & x(101) & x(141) & x(157) & x(160) & x(169) & x(183) & x(186) & x(203) & x(206) & x(207) & x(210) & x(225) & x(227) & x(231) & x(240) & x(255);
    y(212) <= not(p212_out);
    p212 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001100010001110001001101000110",
            TABLE => "111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p212_in,
            y(0) => p212_out,
            y(1 to 14 - 1) => dummy212
        );


    p213_in <= x(5) & x(6) & x(12) & x(19) & x(37) & x(40) & x(45) & x(52) & x(59) & x(62) & x(65) & x(66) & x(76) & x(78) & x(79) & x(82) & x(119) & x(124) & x(126) & x(129) & x(140) & x(143) & x(158) & x(160) & x(214) & x(216) & x(217) & x(245) & x(250) & x(251);
    y(213) <= not(p213_out);
    p213 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011001101000101101111011100000",
            TABLE => "010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p213_in,
            y(0) => p213_out,
            y(1 to 14 - 1) => dummy213
        );


    p214_in <= x(10) & x(21) & x(27) & x(34) & x(50) & x(67) & x(76) & x(82) & x(97) & x(102) & x(110) & x(119) & x(121) & x(133) & x(137) & x(144) & x(152) & x(159) & x(163) & x(165) & x(166) & x(184) & x(189) & x(196) & x(206) & x(208) & x(216) & x(226) & x(233) & x(235) & x(250);
    y(214) <= not(p214_out);
    p214 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111010001010110100001100111011",
            TABLE => "0000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010011101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010010010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101101011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010010000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p214_in,
            y(0) => p214_out,
            y(1 to 14 - 1) => dummy214
        );


    p215_in <= x(7) & x(42) & x(47) & x(69) & x(73) & x(78) & x(80) & x(83) & x(91) & x(118) & x(119) & x(132) & x(134) & x(151) & x(164) & x(219) & x(222) & x(224) & x(234) & x(239) & x(252) & x(253);
    y(215) <= not(p215_out);
    p215 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0101011110101011101111",
            TABLE => "0100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101100000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010010000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p215_in,
            y(0) => p215_out,
            y(1 to 14 - 1) => dummy215
        );


    p216_in <= x(0) & x(1) & x(9) & x(11) & x(25) & x(43) & x(54) & x(64) & x(92) & x(93) & x(97) & x(105) & x(112) & x(113) & x(122) & x(134) & x(139) & x(148) & x(153) & x(169) & x(178) & x(186) & x(196) & x(204) & x(221) & x(222) & x(235) & x(241) & x(242);
    y(216) <= not(p216_out);
    p216 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101001101011011000111101101",
            TABLE => "10110010111110110010000010110010001000001011001000000000001000001011001011011011001001001011001000100100101100100100110100100100100101100110100101101001100101100110100110010110100101100110100100100000101100101011001011111011000000000010000000100000101100100010010010110010101100101101101101001101001001000010010010110010011010011001011010010110011010011001011001101001011010011001011000000010000000000010101100000010001010110000001010111111001010110100001011010100001010110100001000101011010000101011110100101011100101100110100101101001100101100110100110010110100101100110100100010111011111110000000100010111000000010001011100000000000000010001011101111110100000010001011110000001000101111110100010000001100101100110100101101001100101100110100110010110100101100110100101001101110111110000010001001101010011011101101100100100010011010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p216_in,
            y(0) => p216_out,
            y(1 to 13 - 1) => dummy216
        );


    p217_in <= x(13) & x(19) & x(23) & x(24) & x(27) & x(33) & x(35) & x(56) & x(69) & x(78) & x(87) & x(98) & x(112) & x(129) & x(130) & x(135) & x(142) & x(145) & x(146) & x(178) & x(180) & x(201) & x(205) & x(211) & x(217) & x(218) & x(232) & x(238) & x(245) & x(246) & x(252);
    y(217) <= not(p217_out);
    p217 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001011100110111001010010010000",
            TABLE => "1101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010010001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010010000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101101110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p217_in,
            y(0) => p217_out,
            y(1 to 15 - 1) => dummy217
        );


    p218_in <= x(4) & x(14) & x(25) & x(26) & x(28) & x(44) & x(59) & x(62) & x(67) & x(83) & x(87) & x(101) & x(108) & x(112) & x(123) & x(124) & x(149) & x(173) & x(188) & x(206) & x(223) & x(226) & x(234) & x(253);
    y(218) <= not(p218_out);
    p218 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110011010001111011010000",
            TABLE => "000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p218_in,
            y(0) => p218_out,
            y(1 to 14 - 1) => dummy218
        );


    p219_in <= x(47) & x(62) & x(77) & x(88) & x(108) & x(110) & x(135) & x(142) & x(146) & x(155) & x(160) & x(173) & x(179) & x(190) & x(202) & x(222) & x(232) & x(242);
    y(219) <= not(p219_out);
    p219 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010110101101101010",
            TABLE => "001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p219_in,
            y(0) => p219_out,
            y(1 to 14 - 1) => dummy219
        );


    p220_in <= x(10) & x(12) & x(42) & x(46) & x(68) & x(70) & x(81) & x(86) & x(89) & x(91) & x(97) & x(104) & x(108) & x(109) & x(111) & x(116) & x(121) & x(135) & x(137) & x(143) & x(144) & x(156) & x(159) & x(167) & x(178) & x(179) & x(187) & x(205) & x(209) & x(214) & x(216) & x(218) & x(232) & x(233) & x(234) & x(252) & x(255);
    y(220) <= not(p220_out);
    p220 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0101010001001010001001001110001010000",
            TABLE => "0100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101101110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101101000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010011000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101101000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -15,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p220_in,
            y(0) => p220_out,
            y(1 to 15 - 1) => dummy220
        );


    p221_in <= x(34) & x(37) & x(45) & x(50) & x(73) & x(75) & x(81) & x(102) & x(115) & x(129) & x(130) & x(131) & x(140) & x(163) & x(179) & x(188) & x(200) & x(221) & x(226) & x(233) & x(239) & x(249);
    y(221) <= not(p221_out);
    p221 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010111100011001011001",
            TABLE => "0001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010010100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101100100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100100000011010100010000101101010001101001100101100000000000000000",
            SHIFT => 3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p221_in,
            y(0) => p221_out,
            y(1 to 13 - 1) => dummy221
        );


    p222_in <= x(5) & x(16) & x(26) & x(27) & x(34) & x(37) & x(54) & x(68) & x(77) & x(86) & x(101) & x(107) & x(108) & x(111) & x(149) & x(183) & x(188) & x(195) & x(196) & x(197) & x(200) & x(230) & x(242) & x(244) & x(247) & x(250);
    y(222) <= not(p222_out);
    p222 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01011011010111111100000000",
            TABLE => "001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 3,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p222_in,
            y(0) => p222_out,
            y(1 to 13 - 1) => dummy222
        );


    p223_in <= x(9) & x(27) & x(56) & x(57) & x(62) & x(69) & x(77) & x(78) & x(82) & x(119) & x(121) & x(132) & x(134) & x(142) & x(146) & x(160) & x(169) & x(180) & x(182) & x(190) & x(199) & x(202) & x(220) & x(242);
    y(223) <= not(p223_out);
    p223 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010110000101001010100100",
            TABLE => "001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 3,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p223_in,
            y(0) => p223_out,
            y(1 to 13 - 1) => dummy223
        );


    p224_in <= x(25) & x(38) & x(39) & x(47) & x(77) & x(85) & x(90) & x(102) & x(103) & x(114) & x(115) & x(119) & x(129) & x(132) & x(151) & x(156) & x(165) & x(175) & x(188) & x(214) & x(221) & x(232) & x(235) & x(239) & x(251);
    y(224) <= not(p224_out);
    p224 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110111011111001010001111",
            TABLE => "0000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p224_in,
            y(0) => p224_out,
            y(1 to 14 - 1) => dummy224
        );


    p225_in <= x(8) & x(17) & x(25) & x(27) & x(40) & x(42) & x(53) & x(60) & x(62) & x(82) & x(101) & x(113) & x(139) & x(147) & x(153) & x(160) & x(162) & x(165) & x(182) & x(196) & x(205) & x(226) & x(230) & x(231) & x(236) & x(241) & x(251) & x(254);
    y(225) <= not(p225_out);
    p225 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111010111011000111111010010",
            TABLE => "0000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101100000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101101011001000100000101100100010010010010110011010010000000000000000",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p225_in,
            y(0) => p225_out,
            y(1 to 14 - 1) => dummy225
        );


    p226_in <= x(4) & x(25) & x(28) & x(32) & x(57) & x(66) & x(69) & x(76) & x(77) & x(81) & x(85) & x(87) & x(88) & x(93) & x(99) & x(109) & x(124) & x(125) & x(128) & x(154) & x(171) & x(173) & x(180) & x(182) & x(191) & x(198) & x(201) & x(207) & x(209) & x(219) & x(236) & x(237) & x(240) & x(241) & x(242);
    y(226) <= not(p226_out);
    p226 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01010001110100011001101001011001101",
            TABLE => "10001110000010001110111110001110000010000000000010001110000010001000111000011000111001111000111000011000011100011000111000011000100101100110100101101001100101100110100110010110100101100110100100000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100110111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100100100000101100101011001011111011000000000010000000100000101100100010010010110010101100101101101101001101001001000010010010110010011010011001011010010110011010011001011001101001011010011001011000101011000000101011111100101011000000100000000000101011000000100010101101000010101111010010101101000010110101000010101101000010011010011001011010010110011010011001011001101001011010011001011001001101110111110000010001001101010011011101101100100100010011010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 3,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p226_in,
            y(0) => p226_out,
            y(1 to 14 - 1) => dummy226
        );


    p227_in <= x(33) & x(41) & x(49) & x(57) & x(58) & x(74) & x(77) & x(86) & x(87) & x(103) & x(105) & x(120) & x(127) & x(130) & x(134) & x(136) & x(146) & x(172) & x(188) & x(197) & x(199) & x(232);
    y(227) <= not(p227_out);
    p227 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110101010000111000110",
            TABLE => "0000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010011000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p227_in,
            y(0) => p227_out,
            y(1 to 14 - 1) => dummy227
        );


    p228_in <= x(18) & x(26) & x(31) & x(44) & x(50) & x(52) & x(94) & x(112) & x(113) & x(139) & x(154) & x(162) & x(191) & x(203) & x(220) & x(226) & x(227) & x(231) & x(232) & x(234) & x(253);
    y(228) <= not(p228_out);
    p228 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110001100010001110011",
            TABLE => "010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p228_in,
            y(0) => p228_out,
            y(1 to 14 - 1) => dummy228
        );


    p229_in <= x(10) & x(30) & x(50) & x(52) & x(60) & x(66) & x(69) & x(82) & x(97) & x(109) & x(110) & x(112) & x(113) & x(115) & x(123) & x(129) & x(133) & x(139) & x(151) & x(158) & x(186) & x(192) & x(195) & x(196) & x(199) & x(216) & x(226) & x(236) & x(243) & x(246) & x(253);
    y(229) <= not(p229_out);
    p229 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001010000000010101000100111001",
            TABLE => "1101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010011111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010011011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010011011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010010000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 3,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p229_in,
            y(0) => p229_out,
            y(1 to 14 - 1) => dummy229
        );


    p230_in <= x(3) & x(13) & x(41) & x(45) & x(54) & x(61) & x(79) & x(95) & x(104) & x(140) & x(148) & x(164) & x(183) & x(188) & x(196) & x(214) & x(238) & x(241) & x(243) & x(254);
    y(230) <= not(p230_out);
    p230 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000100000100100000",
            TABLE => "110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 4,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p230_in,
            y(0) => p230_out,
            y(1 to 14 - 1) => dummy230
        );


    p231_in <= x(11) & x(15) & x(23) & x(86) & x(92) & x(93) & x(95) & x(96) & x(98) & x(107) & x(121) & x(122) & x(128) & x(133) & x(141) & x(145) & x(146) & x(162) & x(194) & x(197) & x(224) & x(233) & x(245);
    y(231) <= not(p231_out);
    p231 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10100110000111011111101",
            TABLE => "01000000110101000000000001000000110101001111110101000000110101000100001011010100001010110100001011010100101111010100001011010100011010011001011010010110011010011001011001101001011010011001011011010100010000000100000000000000111111011101010011010100010000001101010001000010010000100010101110111101110101001101010001000010100101100110100101101001100101100110100110010110100101100110100100000001000000000001011100000001000101110000000101111111000101111000000111101000000101111000000100010111100000010111111000010111011010011001011010010110011010011001011001101001011010011001011000000100010011010100110111011111001001000100110101001101110110111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p231_in,
            y(0) => p231_out,
            y(1 to 14 - 1) => dummy231
        );


    p232_in <= x(12) & x(16) & x(21) & x(24) & x(36) & x(39) & x(46) & x(48) & x(54) & x(74) & x(99) & x(105) & x(131) & x(142) & x(145) & x(150) & x(167) & x(168) & x(175) & x(187) & x(195) & x(197) & x(209) & x(231) & x(247);
    y(232) <= not(p232_out);
    p232 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111110111011110101001111",
            TABLE => "0000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p232_in,
            y(0) => p232_out,
            y(1 to 14 - 1) => dummy232
        );


    p233_in <= x(12) & x(20) & x(50) & x(52) & x(71) & x(75) & x(80) & x(85) & x(92) & x(98) & x(108) & x(114) & x(119) & x(128) & x(135) & x(145) & x(157) & x(168) & x(185) & x(186) & x(189) & x(194) & x(195) & x(201) & x(202) & x(204) & x(210) & x(219) & x(224) & x(225) & x(237) & x(251);
    y(233) <= not(p233_out);
    p233 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00011111000111110110011010010001",
            TABLE => "011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 3,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p233_in,
            y(0) => p233_out,
            y(1 to 14 - 1) => dummy233
        );


    p234_in <= x(3) & x(6) & x(26) & x(27) & x(44) & x(93) & x(110) & x(129) & x(133) & x(136) & x(139) & x(159) & x(177) & x(181) & x(192) & x(221) & x(226) & x(230) & x(235) & x(236) & x(239) & x(243) & x(247) & x(253);
    y(234) <= not(p234_out);
    p234 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001001001000100110110001",
            TABLE => "110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p234_in,
            y(0) => p234_out,
            y(1 to 13 - 1) => dummy234
        );


    p235_in <= x(16) & x(18) & x(20) & x(24) & x(26) & x(51) & x(55) & x(56) & x(59) & x(62) & x(63) & x(67) & x(69) & x(72) & x(87) & x(106) & x(108) & x(133) & x(144) & x(160) & x(174) & x(186) & x(196) & x(201) & x(206) & x(207) & x(210) & x(227) & x(229) & x(236) & x(240) & x(241) & x(248) & x(249);
    y(235) <= not(p235_out);
    p235 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010110001011101110010011011100101",
            TABLE => "0111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101101101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010010000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101101101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010010000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010100110100000100010011010010010001101001100101100000000000000000",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p235_in,
            y(0) => p235_out,
            y(1 to 15 - 1) => dummy235
        );


    p236_in <= x(12) & x(13) & x(20) & x(28) & x(30) & x(41) & x(46) & x(48) & x(70) & x(73) & x(95) & x(104) & x(111) & x(112) & x(115) & x(127) & x(156) & x(168) & x(176) & x(179) & x(182) & x(189) & x(195) & x(204) & x(215) & x(216) & x(218) & x(231) & x(247) & x(248) & x(254);
    y(236) <= not(p236_out);
    p236 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000111010001000110100101100011",
            TABLE => "0111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101101000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101101011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010010100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => -17,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p236_in,
            y(0) => p236_out,
            y(1 to 15 - 1) => dummy236
        );


    p237_in <= x(4) & x(51) & x(52) & x(66) & x(67) & x(78) & x(79) & x(84) & x(93) & x(95) & x(110) & x(122) & x(128) & x(129) & x(133) & x(140) & x(164) & x(174) & x(201) & x(209) & x(214) & x(217) & x(226) & x(243);
    y(237) <= not(p237_out);
    p237 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000100110010100011001",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p237_in,
            y(0) => p237_out,
            y(1 to 14 - 1) => dummy237
        );


    p238_in <= x(14) & x(15) & x(18) & x(20) & x(22) & x(44) & x(55) & x(67) & x(88) & x(92) & x(98) & x(106) & x(108) & x(111) & x(115) & x(125) & x(127) & x(141) & x(145) & x(153) & x(184) & x(185) & x(189) & x(208) & x(210) & x(213) & x(223) & x(225) & x(227) & x(232) & x(245) & x(248) & x(254);
    y(238) <= not(p238_out);
    p238 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010110011111111111011011110111000",
            TABLE => "001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p238_in,
            y(0) => p238_out,
            y(1 to 14 - 1) => dummy238
        );


    p239_in <= x(1) & x(3) & x(7) & x(11) & x(17) & x(29) & x(34) & x(42) & x(45) & x(58) & x(95) & x(135) & x(143) & x(161) & x(162) & x(164) & x(194) & x(196) & x(236);
    y(239) <= not(p239_out);
    p239 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100100101011101011",
            TABLE => "1011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010010100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101100000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p239_in,
            y(0) => p239_out,
            y(1 to 14 - 1) => dummy239
        );


    p240_in <= x(0) & x(9) & x(33) & x(41) & x(49) & x(65) & x(68) & x(74) & x(76) & x(85) & x(87) & x(101) & x(105) & x(120) & x(121) & x(130) & x(145) & x(150) & x(152) & x(157) & x(174) & x(177) & x(187) & x(188) & x(190) & x(194) & x(198) & x(202) & x(220) & x(229) & x(245) & x(251) & x(252);
    y(240) <= not(p240_out);
    p240 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000000011100110010010111000100100",
            TABLE => "111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110100011101001011011111111",
            SHIFT => 3,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p240_in,
            y(0) => p240_out,
            y(1 to 14 - 1) => dummy240
        );


    p241_in <= x(22) & x(39) & x(45) & x(49) & x(58) & x(60) & x(63) & x(67) & x(77) & x(83) & x(95) & x(103) & x(106) & x(127) & x(138) & x(143) & x(165) & x(183) & x(196) & x(202) & x(213) & x(216) & x(243) & x(250);
    y(241) <= not(p241_out);
    p241 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010110101001001100110101",
            TABLE => "001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p241_in,
            y(0) => p241_out,
            y(1 to 14 - 1) => dummy241
        );


    p242_in <= x(27) & x(30) & x(55) & x(62) & x(67) & x(79) & x(87) & x(91) & x(110) & x(112) & x(124) & x(136) & x(142) & x(154) & x(181) & x(190) & x(198) & x(218) & x(238) & x(246) & x(247);
    y(242) <= not(p242_out);
    p242 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101101001101101101111",
            TABLE => "000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p242_in,
            y(0) => p242_out,
            y(1 to 14 - 1) => dummy242
        );


    p243_in <= x(43) & x(57) & x(59) & x(76) & x(83) & x(85) & x(101) & x(130) & x(141) & x(145) & x(188) & x(193) & x(207) & x(236) & x(247);
    y(243) <= not(p243_out);
    p243 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100001110100011",
            TABLE => "110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p243_in,
            y(0) => p243_out,
            y(1 to 13 - 1) => dummy243
        );


    p244_in <= x(14) & x(15) & x(22) & x(24) & x(33) & x(36) & x(44) & x(55) & x(58) & x(61) & x(67) & x(69) & x(78) & x(79) & x(97) & x(113) & x(117) & x(123) & x(124) & x(127) & x(131) & x(141) & x(145) & x(155) & x(165) & x(167) & x(174) & x(187) & x(191) & x(198) & x(199) & x(213);
    y(244) <= not(p244_out);
    p244 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10010111100001001100101100010000",
            TABLE => "010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 3,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p244_in,
            y(0) => p244_out,
            y(1 to 14 - 1) => dummy244
        );


    p245_in <= x(22) & x(23) & x(27) & x(33) & x(35) & x(36) & x(60) & x(72) & x(78) & x(98) & x(99) & x(111) & x(119) & x(124) & x(135) & x(142) & x(145) & x(181) & x(182) & x(198) & x(210) & x(213) & x(217) & x(218) & x(221) & x(225) & x(232) & x(237) & x(245);
    y(245) <= not(p245_out);
    p245 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01100101101010011110001100001",
            TABLE => "01000000110101001101010011111101000000000100000001000000110101000100001011010100110101001011110100101011010000100100001011010100011010011001011010010110011010011001011001101001011010011001011000100000101100101011001011111011000000000010000000100000101100100010010010110010101100101101101101001101001001000010010010110010011010011001011010010110011010011001011001101001011010011001011000010111000000010000000100000000011111110001011100010111000000010001011110000001100000011110100001111110000101110001011110000001100101100110100101101001100101100110100110010110100101100110100101110001000100000001000000000000111101110111000101110001000100000111000100011000000110001000111011100111011100010111000100011000011010011001011010010110011010011001011001101001011010011001011011111101110101001101010001000000101111011101010011010100010000100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p245_in,
            y(0) => p245_out,
            y(1 to 14 - 1) => dummy245
        );


    p246_in <= x(25) & x(44) & x(52) & x(67) & x(79) & x(80) & x(84) & x(95) & x(108) & x(111) & x(114) & x(135) & x(136) & x(140) & x(149) & x(164) & x(178) & x(181) & x(196) & x(214) & x(217) & x(243) & x(253) & x(254);
    y(246) <= not(p246_out);
    p246 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101101100011000100101010",
            TABLE => "000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 3,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p246_in,
            y(0) => p246_out,
            y(1 to 13 - 1) => dummy246
        );


    p247_in <= x(2) & x(6) & x(9) & x(12) & x(18) & x(28) & x(38) & x(44) & x(51) & x(52) & x(68) & x(69) & x(92) & x(102) & x(108) & x(125) & x(134) & x(147) & x(154) & x(156) & x(173) & x(179) & x(184) & x(191) & x(193) & x(197) & x(205) & x(211) & x(230) & x(232) & x(251);
    y(247) <= not(p247_out);
    p247 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100101101100000011000000110001",
            TABLE => "0010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101100000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101101110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101101000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 3,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p247_in,
            y(0) => p247_out,
            y(1 to 14 - 1) => dummy247
        );


    p248_in <= x(4) & x(6) & x(19) & x(20) & x(23) & x(33) & x(35) & x(40) & x(52) & x(54) & x(66) & x(76) & x(87) & x(119) & x(127) & x(131) & x(142) & x(166) & x(175) & x(177) & x(179) & x(182) & x(192) & x(212) & x(218) & x(222) & x(248) & x(250);
    y(248) <= not(p248_out);
    p248 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0101011101011010010010110010",
            TABLE => "0100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101100000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101101011001000100000101100100010010010010110011010010000000000000000",
            SHIFT => 4,
            B => -12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p248_in,
            y(0) => p248_out,
            y(1 to 14 - 1) => dummy248
        );


    p249_in <= x(17) & x(25) & x(27) & x(33) & x(52) & x(59) & x(62) & x(68) & x(83) & x(86) & x(94) & x(104) & x(119) & x(138) & x(148) & x(151) & x(156) & x(160) & x(166) & x(168) & x(171) & x(176) & x(177) & x(195) & x(203) & x(205) & x(215) & x(217) & x(240) & x(247);
    y(249) <= not(p249_out);
    p249 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010001000000000111001110100111",
            TABLE => "110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p249_in,
            y(0) => p249_out,
            y(1 to 15 - 1) => dummy249
        );


    p250_in <= x(8) & x(18) & x(28) & x(29) & x(31) & x(49) & x(51) & x(68) & x(84) & x(89) & x(90) & x(91) & x(104) & x(125) & x(126) & x(155) & x(156) & x(162) & x(177) & x(179) & x(191) & x(201) & x(205) & x(213) & x(217) & x(226);
    y(250) <= not(p250_out);
    p250 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11000101010000000000001000",
            TABLE => "010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 3,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p250_in,
            y(0) => p250_out,
            y(1 to 13 - 1) => dummy250
        );


    p251_in <= x(9) & x(12) & x(28) & x(30) & x(36) & x(43) & x(44) & x(49) & x(67) & x(73) & x(82) & x(100) & x(134) & x(141) & x(145) & x(146) & x(147) & x(180) & x(199) & x(202) & x(211) & x(212) & x(255);
    y(251) <= not(p251_out);
    p251 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101110010100111001011",
            TABLE => "01110001111101110001000001110001000100000111000100000000000100000111000111100111000110000111000100011000011100011000111000011000011010011001011010010110011010011001011001101001011010011001011001001101000001000000010000000000110111110100110101001101000001000100110100100100001001001011001011011011010011010100110100100100011010011001011010010110011010011001011001101001011010011001011000101011101111110000001000101011000000100010101100000000000000100010101110111101010000100010101101000010001010111101010001000010011010011001011010010110011010011001011001101001011010011001011001110001111101110001000001110001011100011110011100011000011100010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 3,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p251_in,
            y(0) => p251_out,
            y(1 to 13 - 1) => dummy251
        );


    p252_in <= x(12) & x(16) & x(18) & x(26) & x(46) & x(63) & x(67) & x(98) & x(104) & x(105) & x(108) & x(117) & x(137) & x(142) & x(146) & x(153) & x(158) & x(167) & x(170) & x(175) & x(179) & x(181) & x(182) & x(205) & x(212) & x(224) & x(234) & x(248) & x(252);
    y(252) <= not(p252_out);
    p252 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110100110001001111011100101",
            TABLE => "00000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100110001110111011110000100010001110000010001000111000000000000010001000111011100111000110001000111000011000100011100111000100011000100101100110100101101001100101100110100110010110100101100110100101110001000100001111011101110001000100000000000001110001000100000111000100011000111001110111000100011000100011100111000100011000011010011001011010010110011010011001011001101001011010011001011000000001000000000001011100000001000101110000000101111111000101111000000111101000000101111000000100010111100000010111111000010111011010011001011010010110011010011001011001101001011010011001011011011111010011010100110100000100110110110100110101001101001001001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p252_in,
            y(0) => p252_out,
            y(1 to 14 - 1) => dummy252
        );


    p253_in <= x(9) & x(14) & x(46) & x(50) & x(70) & x(74) & x(77) & x(78) & x(86) & x(90) & x(96) & x(101) & x(105) & x(107) & x(111) & x(112) & x(130) & x(132) & x(134) & x(142) & x(146) & x(151) & x(153) & x(154) & x(188) & x(212) & x(222) & x(231) & x(252);
    y(253) <= not(p253_out);
    p253 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101100101011100100111111000",
            TABLE => "01110001111101110001000001110001000100000111000100000000000100000111000111100111000110000111000100011000011100011000111000011000011010011001011010010110011010011001011001101001011010011001011010110010111110110010000010110010001000001011001000000000001000001011001011011011001001001011001000100100101100100100110100100100100101100110100101101001100101100110100110010110100101100110100100000000010000000100000011010100010000001101010011010100111111010010101101000010010000101101010001000010110101001101010010111101100101100110100101101001100101100110100110010110100101100110100100010111011111110000000100010111000000010001011100000000000000010001011101111110100000010001011110000001000101111110100010000001100101100110100101101001100101100110100110010110100101100110100110000000111010001110100011111110100000011110100011101000011111101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 3,
            B => -11,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p253_in,
            y(0) => p253_out,
            y(1 to 13 - 1) => dummy253
        );


    p254_in <= x(7) & x(8) & x(13) & x(28) & x(40) & x(59) & x(70) & x(88) & x(91) & x(101) & x(130) & x(134) & x(147) & x(160) & x(166) & x(168) & x(173) & x(176) & x(183) & x(186) & x(189) & x(190) & x(199) & x(216) & x(223) & x(228) & x(230) & x(254);
    y(254) <= not(p254_out);
    p254 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100111000001111000001111011",
            TABLE => "0001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010011110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101100000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100001000001110001000110000111000110010110011010010000000000000000",
            SHIFT => 3,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p254_in,
            y(0) => p254_out,
            y(1 to 13 - 1) => dummy254
        );


    p255_in <= x(10) & x(32) & x(52) & x(54) & x(60) & x(66) & x(81) & x(82) & x(95) & x(97) & x(102) & x(113) & x(122) & x(156) & x(176) & x(184) & x(186) & x(195) & x(197) & x(203) & x(204) & x(205) & x(209) & x(214) & x(216) & x(219) & x(242);
    y(255) <= not(p255_out);
    p255 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110110111101001010111111001",
            TABLE => "000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001110101001001011011111111",
            SHIFT => 3,
            B => 12,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p255_in,
            y(0) => p255_out,
            y(1 to 13 - 1) => dummy255
        );



end layer_3;

architecture layer_4 of layer is

    Component perceptron
    Generic (
        WEIGHTS : STD_LOGIC_VECTOR;
        SHIFT : Integer;     -- number of shift (left + or right -)
        B : Integer;          -- bias of batch norm
        BATCH_POSITIVE : Boolean    
    );
    Port ( 
        x : in STD_LOGIC_VECTOR;
        y : out STD_LOGIC_VECTOR
   );
    end component;
    
    -- Signals
    signal p0_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p0_out : STD_LOGIC;
	signal p1_in : STD_LOGIC_VECTOR(0 to 14 - 1);
	signal p1_out : STD_LOGIC;
	signal p2_in : STD_LOGIC_VECTOR(0 to 12 - 1);
	signal p2_out : STD_LOGIC;
	signal p3_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p3_out : STD_LOGIC;
	signal p4_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p4_out : STD_LOGIC;
	signal p5_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p5_out : STD_LOGIC;
	signal p6_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p6_out : STD_LOGIC;
	signal p7_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p7_out : STD_LOGIC;
	signal p8_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p8_out : STD_LOGIC;
	signal p9_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p9_out : STD_LOGIC;
	signal p10_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p10_out : STD_LOGIC;
	signal p11_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p11_out : STD_LOGIC;
	signal p12_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p12_out : STD_LOGIC;
	signal p13_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p13_out : STD_LOGIC;
	signal p14_in : STD_LOGIC_VECTOR(0 to 11 - 1);
	signal p14_out : STD_LOGIC;
	signal p15_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p15_out : STD_LOGIC;
	signal p16_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p16_out : STD_LOGIC;
	signal p17_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p17_out : STD_LOGIC;
	signal p18_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p18_out : STD_LOGIC;
	signal p19_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p19_out : STD_LOGIC;
	signal p20_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p20_out : STD_LOGIC;
	signal p21_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p21_out : STD_LOGIC;
	signal p22_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p22_out : STD_LOGIC;
	signal p23_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p23_out : STD_LOGIC;
	signal p24_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p24_out : STD_LOGIC;
	signal p25_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p25_out : STD_LOGIC;
	signal p26_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p26_out : STD_LOGIC;
	signal p27_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p27_out : STD_LOGIC;
	signal p28_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p28_out : STD_LOGIC;
	signal p29_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p29_out : STD_LOGIC;
	signal p30_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p30_out : STD_LOGIC;
	signal p31_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p31_out : STD_LOGIC;
	signal p32_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p32_out : STD_LOGIC;
	signal p33_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p33_out : STD_LOGIC;
	signal p34_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p34_out : STD_LOGIC;
	signal p35_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p35_out : STD_LOGIC;
	signal p36_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p36_out : STD_LOGIC;
	signal p37_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p37_out : STD_LOGIC;
	signal p38_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p38_out : STD_LOGIC;
	signal p39_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p39_out : STD_LOGIC;
	signal p40_in : STD_LOGIC_VECTOR(0 to 13 - 1);
	signal p40_out : STD_LOGIC;
	signal p41_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p41_out : STD_LOGIC;
	signal p42_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p42_out : STD_LOGIC;
	signal p43_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p43_out : STD_LOGIC;
	signal p44_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p44_out : STD_LOGIC;
	signal p45_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p45_out : STD_LOGIC;
	signal p46_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p46_out : STD_LOGIC;
	signal p47_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p47_out : STD_LOGIC;
	signal p48_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p48_out : STD_LOGIC;
	signal p49_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p49_out : STD_LOGIC;
	signal p50_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p50_out : STD_LOGIC;
	signal p51_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p51_out : STD_LOGIC;
	signal p52_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p52_out : STD_LOGIC;
	signal p53_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p53_out : STD_LOGIC;
	signal p54_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p54_out : STD_LOGIC;
	signal p55_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p55_out : STD_LOGIC;
	signal p56_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p56_out : STD_LOGIC;
	signal p57_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p57_out : STD_LOGIC;
	signal p58_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p58_out : STD_LOGIC;
	signal p59_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p59_out : STD_LOGIC;
	signal p60_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p60_out : STD_LOGIC;
	signal p62_in : STD_LOGIC_VECTOR(0 to 14 - 1);
	signal p62_out : STD_LOGIC;
	signal p63_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p63_out : STD_LOGIC;
	signal p64_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p64_out : STD_LOGIC;
	signal p65_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p65_out : STD_LOGIC;
	signal p66_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p66_out : STD_LOGIC;
	signal p67_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p67_out : STD_LOGIC;
	signal p68_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p68_out : STD_LOGIC;
	signal p69_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p69_out : STD_LOGIC;
	signal p70_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p70_out : STD_LOGIC;
	signal p71_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p71_out : STD_LOGIC;
	signal p72_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p72_out : STD_LOGIC;
	signal p73_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p73_out : STD_LOGIC;
	signal p74_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p74_out : STD_LOGIC;
	signal p75_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p75_out : STD_LOGIC;
	signal p76_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p76_out : STD_LOGIC;
	signal p77_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p77_out : STD_LOGIC;
	signal p78_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p78_out : STD_LOGIC;
	signal p79_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p79_out : STD_LOGIC;
	signal p80_in : STD_LOGIC_VECTOR(0 to 14 - 1);
	signal p80_out : STD_LOGIC;
	signal p81_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p81_out : STD_LOGIC;
	signal p82_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p82_out : STD_LOGIC;
	signal p83_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p83_out : STD_LOGIC;
	signal p84_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p84_out : STD_LOGIC;
	signal p85_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p85_out : STD_LOGIC;
	signal p86_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p86_out : STD_LOGIC;
	signal p87_in : STD_LOGIC_VECTOR(0 to 29 - 1);
	signal p87_out : STD_LOGIC;
	signal p88_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p88_out : STD_LOGIC;
	signal p89_in : STD_LOGIC_VECTOR(0 to 35 - 1);
	signal p89_out : STD_LOGIC;
	signal p90_in : STD_LOGIC_VECTOR(0 to 6 - 1);
	signal p90_out : STD_LOGIC;
	signal p91_in : STD_LOGIC_VECTOR(0 to 14 - 1);
	signal p91_out : STD_LOGIC;
	signal p92_in : STD_LOGIC_VECTOR(0 to 13 - 1);
	signal p92_out : STD_LOGIC;
	signal p93_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p93_out : STD_LOGIC;
	signal p94_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p94_out : STD_LOGIC;
	signal p95_in : STD_LOGIC_VECTOR(0 to 14 - 1);
	signal p95_out : STD_LOGIC;
	signal p96_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p96_out : STD_LOGIC;
	signal p97_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p97_out : STD_LOGIC;
	signal p98_in : STD_LOGIC_VECTOR(0 to 4 - 1);
	signal p98_out : STD_LOGIC;
	signal p99_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p99_out : STD_LOGIC;
	signal p100_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p100_out : STD_LOGIC;
	signal p101_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p101_out : STD_LOGIC;
	signal p102_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p102_out : STD_LOGIC;
	signal p103_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p103_out : STD_LOGIC;
	signal p104_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p104_out : STD_LOGIC;
	signal p105_in : STD_LOGIC_VECTOR(0 to 12 - 1);
	signal p105_out : STD_LOGIC;
	signal p106_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p106_out : STD_LOGIC;
	signal p107_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p107_out : STD_LOGIC;
	signal p108_in : STD_LOGIC_VECTOR(0 to 14 - 1);
	signal p108_out : STD_LOGIC;
	signal p109_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p109_out : STD_LOGIC;
	signal p110_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p110_out : STD_LOGIC;
	signal p111_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p111_out : STD_LOGIC;
	signal p112_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p112_out : STD_LOGIC;
	signal p113_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p113_out : STD_LOGIC;
	signal p114_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p114_out : STD_LOGIC;
	signal p115_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p115_out : STD_LOGIC;
	signal p116_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p116_out : STD_LOGIC;
	signal p117_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p117_out : STD_LOGIC;
	signal p118_in : STD_LOGIC_VECTOR(0 to 13 - 1);
	signal p118_out : STD_LOGIC;
	signal p119_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p119_out : STD_LOGIC;
	signal p120_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p120_out : STD_LOGIC;
	signal p121_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p121_out : STD_LOGIC;
	signal p122_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p122_out : STD_LOGIC;
	signal p123_in : STD_LOGIC_VECTOR(0 to 12 - 1);
	signal p123_out : STD_LOGIC;
	signal p124_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p124_out : STD_LOGIC;
	signal p125_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p125_out : STD_LOGIC;
	signal p126_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p126_out : STD_LOGIC;
	signal p127_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p127_out : STD_LOGIC;
	signal p128_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p128_out : STD_LOGIC;
	signal p129_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p129_out : STD_LOGIC;
	signal p130_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p130_out : STD_LOGIC;
	signal p131_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p131_out : STD_LOGIC;
	signal p132_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p132_out : STD_LOGIC;
	signal p133_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p133_out : STD_LOGIC;
	signal p134_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p134_out : STD_LOGIC;
	signal p135_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p135_out : STD_LOGIC;
	signal p136_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p136_out : STD_LOGIC;
	signal p137_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p137_out : STD_LOGIC;
	signal p138_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p138_out : STD_LOGIC;
	signal p139_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p139_out : STD_LOGIC;
	signal p140_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p140_out : STD_LOGIC;
	signal p141_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p141_out : STD_LOGIC;
	signal p142_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p142_out : STD_LOGIC;
	signal p143_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p143_out : STD_LOGIC;
	signal p144_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p144_out : STD_LOGIC;
	signal p145_in : STD_LOGIC_VECTOR(0 to 13 - 1);
	signal p145_out : STD_LOGIC;
	signal p146_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p146_out : STD_LOGIC;
	signal p147_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p147_out : STD_LOGIC;
	signal p148_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p148_out : STD_LOGIC;
	signal p149_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p149_out : STD_LOGIC;
	signal p150_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p150_out : STD_LOGIC;
	signal p151_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p151_out : STD_LOGIC;
	signal p152_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p152_out : STD_LOGIC;
	signal p153_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p153_out : STD_LOGIC;
	signal p154_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p154_out : STD_LOGIC;
	signal p155_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p155_out : STD_LOGIC;
	signal p156_in : STD_LOGIC_VECTOR(0 to 10 - 1);
	signal p156_out : STD_LOGIC;
	signal p157_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p157_out : STD_LOGIC;
	signal p158_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p158_out : STD_LOGIC;
	signal p159_in : STD_LOGIC_VECTOR(0 to 31 - 1);
	signal p159_out : STD_LOGIC;
	signal p160_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p160_out : STD_LOGIC;
	signal p161_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p161_out : STD_LOGIC;
	signal p162_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p162_out : STD_LOGIC;
	signal p163_in : STD_LOGIC_VECTOR(0 to 11 - 1);
	signal p163_out : STD_LOGIC;
	signal p164_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p164_out : STD_LOGIC;
	signal p165_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p165_out : STD_LOGIC;
	signal p166_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p166_out : STD_LOGIC;
	signal p167_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p167_out : STD_LOGIC;
	signal p168_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p168_out : STD_LOGIC;
	signal p169_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p169_out : STD_LOGIC;
	signal p170_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p170_out : STD_LOGIC;
	signal p171_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p171_out : STD_LOGIC;
	signal p172_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p172_out : STD_LOGIC;
	signal p173_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p173_out : STD_LOGIC;
	signal p174_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p174_out : STD_LOGIC;
	signal p175_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p175_out : STD_LOGIC;
	signal p176_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p176_out : STD_LOGIC;
	signal p177_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p177_out : STD_LOGIC;
	signal p178_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p178_out : STD_LOGIC;
	signal p179_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p179_out : STD_LOGIC;
	signal p180_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p180_out : STD_LOGIC;
	signal p181_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p181_out : STD_LOGIC;
	signal p182_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p182_out : STD_LOGIC;
	signal p183_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p183_out : STD_LOGIC;
	signal p184_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p184_out : STD_LOGIC;
	signal p185_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p185_out : STD_LOGIC;
	signal p186_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p186_out : STD_LOGIC;
	signal p187_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p187_out : STD_LOGIC;
	signal p188_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p188_out : STD_LOGIC;
	signal p189_in : STD_LOGIC_VECTOR(0 to 14 - 1);
	signal p189_out : STD_LOGIC;
	signal p190_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p190_out : STD_LOGIC;
	signal p191_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p191_out : STD_LOGIC;
	signal p192_in : STD_LOGIC_VECTOR(0 to 14 - 1);
	signal p192_out : STD_LOGIC;
	signal p193_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p193_out : STD_LOGIC;
	signal p194_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p194_out : STD_LOGIC;
	signal p195_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p195_out : STD_LOGIC;
	signal p196_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p196_out : STD_LOGIC;
	signal p197_in : STD_LOGIC_VECTOR(0 to 5 - 1);
	signal p197_out : STD_LOGIC;
	signal p198_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p198_out : STD_LOGIC;
	signal p199_in : STD_LOGIC_VECTOR(0 to 33 - 1);
	signal p199_out : STD_LOGIC;
	signal p200_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p200_out : STD_LOGIC;
	signal p201_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p201_out : STD_LOGIC;
	signal p202_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p202_out : STD_LOGIC;
	signal p203_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p203_out : STD_LOGIC;
	signal p204_in : STD_LOGIC_VECTOR(0 to 8 - 1);
	signal p204_out : STD_LOGIC;
	signal p205_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p205_out : STD_LOGIC;
	signal p206_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p206_out : STD_LOGIC;
	signal p207_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p207_out : STD_LOGIC;
	signal p208_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p208_out : STD_LOGIC;
	signal p209_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p209_out : STD_LOGIC;
	signal p210_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p210_out : STD_LOGIC;
	signal p211_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p211_out : STD_LOGIC;
	signal p212_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p212_out : STD_LOGIC;
	signal p213_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p213_out : STD_LOGIC;
	signal p214_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p214_out : STD_LOGIC;
	signal p215_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p215_out : STD_LOGIC;
	signal p216_in : STD_LOGIC_VECTOR(0 to 9 - 1);
	signal p216_out : STD_LOGIC;
	signal p217_in : STD_LOGIC_VECTOR(0 to 26 - 1);
	signal p217_out : STD_LOGIC;
	signal p218_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p218_out : STD_LOGIC;
	signal p219_in : STD_LOGIC_VECTOR(0 to 28 - 1);
	signal p219_out : STD_LOGIC;
	signal p220_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p220_out : STD_LOGIC;
	signal p221_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p221_out : STD_LOGIC;
	signal p222_in : STD_LOGIC_VECTOR(0 to 21 - 1);
	signal p222_out : STD_LOGIC;
	signal p223_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p223_out : STD_LOGIC;
	signal p224_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p224_out : STD_LOGIC;
	signal p225_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p225_out : STD_LOGIC;
	signal p226_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p226_out : STD_LOGIC;
	signal p227_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p227_out : STD_LOGIC;
	signal p228_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p228_out : STD_LOGIC;
	signal p229_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p229_out : STD_LOGIC;
	signal p230_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p230_out : STD_LOGIC;
	signal p231_in : STD_LOGIC_VECTOR(0 to 15 - 1);
	signal p231_out : STD_LOGIC;
	signal p232_in : STD_LOGIC_VECTOR(0 to 7 - 1);
	signal p232_out : STD_LOGIC;
	signal p233_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p233_out : STD_LOGIC;
	signal p234_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p234_out : STD_LOGIC;
	signal p235_in : STD_LOGIC_VECTOR(0 to 22 - 1);
	signal p235_out : STD_LOGIC;
	signal p236_in : STD_LOGIC_VECTOR(0 to 17 - 1);
	signal p236_out : STD_LOGIC;
	signal p237_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p237_out : STD_LOGIC;
	signal p238_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p238_out : STD_LOGIC;
	signal p239_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p239_out : STD_LOGIC;
	signal p240_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p240_out : STD_LOGIC;
	signal p241_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p241_out : STD_LOGIC;
	signal p242_in : STD_LOGIC_VECTOR(0 to 20 - 1);
	signal p242_out : STD_LOGIC;
	signal p243_in : STD_LOGIC_VECTOR(0 to 14 - 1);
	signal p243_out : STD_LOGIC;
	signal p244_in : STD_LOGIC_VECTOR(0 to 24 - 1);
	signal p244_out : STD_LOGIC;
	signal p245_in : STD_LOGIC_VECTOR(0 to 23 - 1);
	signal p245_out : STD_LOGIC;
	signal p246_in : STD_LOGIC_VECTOR(0 to 32 - 1);
	signal p246_out : STD_LOGIC;
	signal p247_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p247_out : STD_LOGIC;
	signal p248_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p248_out : STD_LOGIC;
	signal p249_in : STD_LOGIC_VECTOR(0 to 16 - 1);
	signal p249_out : STD_LOGIC;
	signal p250_in : STD_LOGIC_VECTOR(0 to 18 - 1);
	signal p250_out : STD_LOGIC;
	signal p251_in : STD_LOGIC_VECTOR(0 to 25 - 1);
	signal p251_out : STD_LOGIC;
	signal p252_in : STD_LOGIC_VECTOR(0 to 27 - 1);
	signal p252_out : STD_LOGIC;
	signal p253_in : STD_LOGIC_VECTOR(0 to 30 - 1);
	signal p253_out : STD_LOGIC;
	signal p254_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p254_out : STD_LOGIC;
	signal p255_in : STD_LOGIC_VECTOR(0 to 19 - 1);
	signal p255_out : STD_LOGIC;
	
    
    -- Dummies
    signal dummy0 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy1 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy2 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy3 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy4 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy5 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy6 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy7 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy8 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy9 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy10 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy11 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy12 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy13 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy14 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy15 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy16 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy17 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy18 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy19 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy20 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy21 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy22 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy23 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy24 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy25 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy26 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy27 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy28 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy29 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy30 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy31 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy32 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy33 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy34 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy35 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy36 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy37 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy38 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy39 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy40 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy41 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy42 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy43 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy44 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy45 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy46 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy47 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy48 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy49 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy50 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy51 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy52 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy53 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy54 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy55 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy56 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy57 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy58 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy59 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy60 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy62 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy63 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy64 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy65 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy66 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy67 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy68 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy69 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy70 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy71 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy72 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy73 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy74 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy75 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy76 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy77 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy78 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy79 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy80 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy81 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy82 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy83 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy84 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy85 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy86 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy87 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy88 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy89 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy90 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy91 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy92 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy93 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy94 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy95 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy96 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy97 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy98 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy99 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy100 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy101 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy102 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy103 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy104 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy105 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy106 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy107 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy108 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy109 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy110 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy111 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy112 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy113 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy114 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy115 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy116 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy117 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy118 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy119 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy120 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy121 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy122 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy123 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy124 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy125 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy126 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy127 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy128 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy129 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy130 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy131 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy132 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy133 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy134 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy135 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy136 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy137 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy138 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy139 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy140 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy141 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy142 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy143 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy144 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy145 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy146 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy147 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy148 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy149 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy150 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy151 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy152 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy153 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy154 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy155 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy156 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy157 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy158 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy159 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy160 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy161 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy162 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy163 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy164 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy165 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy166 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy167 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy168 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy169 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy170 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy171 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy172 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy173 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy174 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy175 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy176 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy177 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy178 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy179 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy180 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy181 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy182 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy183 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy184 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy185 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy186 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy187 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy188 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy189 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy190 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy191 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy192 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy193 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy194 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy195 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy196 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy197 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy198 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy199 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy200 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy201 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy202 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy203 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy204 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy205 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy206 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy207 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy208 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy209 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy210 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy211 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy212 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy213 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy214 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy215 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy216 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy217 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy218 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy219 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy220 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy221 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy222 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy223 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy224 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy225 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy226 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy227 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy228 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy229 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy230 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy231 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy232 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy233 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy234 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy235 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy236 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy237 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy238 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy239 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy240 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy241 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy242 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy243 : STD_LOGIC_VECTOR(0 to 13 - 2);
	signal dummy244 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy245 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy246 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy247 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy248 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy249 : STD_LOGIC_VECTOR(0 to 15 - 2);
	signal dummy250 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy251 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy252 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy253 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy254 : STD_LOGIC_VECTOR(0 to 14 - 2);
	signal dummy255 : STD_LOGIC_VECTOR(0 to 14 - 2);
	 

begin

    
    p0_in <= x(17) & x(27) & x(36) & x(40) & x(49) & x(51) & x(56) & x(68) & x(78) & x(80) & x(97) & x(100) & x(103) & x(128) & x(131) & x(135) & x(137) & x(138) & x(145) & x(148) & x(172) & x(177) & x(178) & x(222) & x(223) & x(227) & x(240) & x(251) & x(252) & x(253) & x(254);
    y(0) <= not(p0_out);
    p0 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001011101000000010111011011010",
            TABLE => "0100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101101111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p0_in,
            y(0) => p0_out,
            y(1 to 15 - 1) => dummy0
        );


    p1_in <= x(11) & x(16) & x(48) & x(49) & x(51) & x(65) & x(91) & x(101) & x(111) & x(174) & x(187) & x(198) & x(213) & x(239);
    y(1) <= not(p1_out);
    p1 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000011001110",
            TABLE => "111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p1_in,
            y(0) => p1_out,
            y(1 to 14 - 1) => dummy1
        );


    p2_in <= x(35) & x(38) & x(47) & x(85) & x(121) & x(152) & x(183) & x(191) & x(203) & x(206) & x(226) & x(249);
    y(2) <= not(p2_out);
    p2 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100100010011",
            TABLE => "100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p2_in,
            y(0) => p2_out,
            y(1 to 13 - 1) => dummy2
        );


    p3_in <= x(5) & x(18) & x(21) & x(32) & x(37) & x(52) & x(62) & x(89) & x(98) & x(102) & x(105) & x(107) & x(126) & x(130) & x(173) & x(208) & x(216) & x(221) & x(224) & x(234) & x(239) & x(251);
    y(3) <= not(p3_out);
    p3 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0011100100111101101010",
            TABLE => "0010101110111111000000100010101100000010001010110000000000000010001010111011110101000010001010110100001000101011110101000100001001101001100101101001011001101001100101100110100101101001100101100111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101100000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010010010000010110010001001001011001001101001100101100000000000000000",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p3_in,
            y(0) => p3_out,
            y(1 to 14 - 1) => dummy3
        );


    p4_in <= x(4) & x(10) & x(15) & x(18) & x(24) & x(26) & x(44) & x(69) & x(89) & x(110) & x(144) & x(146) & x(162) & x(170) & x(192) & x(213) & x(241);
    y(4) <= not(p4_out);
    p4 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00010110101100010",
            TABLE => "11011111010011010100110100000100010011010000010000000100000000001101101101001101010011010010010001001101001001000010010010110010100101100110100101101001100101100110100110010110100101100110100100010000011100010000000000010000011100011111011100010000011100010001100001110001100011100001100001110001111001110001100001110001100101100110100101101001100101100110100110010110100101100110100111111011101100101011001000100000110110111011001010110010001001000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p4_in,
            y(0) => p4_out,
            y(1 to 14 - 1) => dummy4
        );


    p5_in <= x(6) & x(29) & x(55) & x(56) & x(75) & x(88) & x(93) & x(105) & x(112) & x(117) & x(141) & x(152) & x(174) & x(198) & x(200) & x(204) & x(218) & x(228) & x(237) & x(253);
    y(5) <= not(p5_out);
    p5 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01011001100101001010",
            TABLE => "001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p5_in,
            y(0) => p5_out,
            y(1 to 14 - 1) => dummy5
        );


    p6_in <= x(16) & x(31) & x(34) & x(43) & x(49) & x(59) & x(65) & x(89) & x(92) & x(103) & x(120) & x(121) & x(123) & x(125) & x(138) & x(147) & x(153) & x(158) & x(171) & x(185) & x(205) & x(212) & x(253);
    y(6) <= not(p6_out);
    p6 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00000100110101111110010",
            TABLE => "11111101110101001101010001000000110101000100000001000000000000001011110111010100110101000100001011010100010000100100001000101011011010011001011010010110011010011001011001101001011010011001011001001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011000000001000101110001011101111111000000000000000100000001000101111000000100010111000101110111111011101000100000011000000100010111011010011001011010010110011010011001011001101001011010011001011010110010001000001111101110110010101100100010010011011011101100101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p6_in,
            y(0) => p6_out,
            y(1 to 14 - 1) => dummy6
        );


    p7_in <= x(11) & x(14) & x(22) & x(32) & x(35) & x(40) & x(47) & x(48) & x(51) & x(54) & x(62) & x(70) & x(74) & x(84) & x(87) & x(91) & x(97) & x(117) & x(125) & x(132) & x(140) & x(141) & x(143) & x(196) & x(215) & x(230) & x(239) & x(240) & x(244) & x(246);
    y(7) <= not(p7_out);
    p7 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001100110101100011000110111001",
            TABLE => "100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p7_in,
            y(0) => p7_out,
            y(1 to 14 - 1) => dummy7
        );


    p8_in <= x(9) & x(27) & x(178) & x(186) & x(198);
    y(8) <= not(p8_out);
    p8 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11110",
            TABLE => "00000010001010110010101110111111010000100010101100101011101111011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p8_in,
            y(0) => p8_out,
            y(1 to 13 - 1) => dummy8
        );


    p9_in <= x(0) & x(8) & x(17) & x(30) & x(31) & x(54) & x(70) & x(71) & x(78) & x(80) & x(91) & x(95) & x(97) & x(103) & x(118) & x(121) & x(123) & x(125) & x(132) & x(138) & x(141) & x(143) & x(160) & x(164) & x(180) & x(183) & x(201) & x(210) & x(236) & x(238) & x(239) & x(244);
    y(9) <= not(p9_out);
    p9 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10110000011101110111000101101001",
            TABLE => "000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p9_in,
            y(0) => p9_out,
            y(1 to 15 - 1) => dummy9
        );


    p10_in <= x(5) & x(11) & x(14) & x(28) & x(29) & x(40) & x(41) & x(47) & x(50) & x(51) & x(70) & x(88) & x(89) & x(104) & x(126) & x(131) & x(140) & x(142) & x(179) & x(186) & x(196) & x(232) & x(240) & x(255);
    y(10) <= not(p10_out);
    p10 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011111000100111010001111",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p10_in,
            y(0) => p10_out,
            y(1 to 14 - 1) => dummy10
        );


    p11_in <= x(14) & x(16) & x(37) & x(48) & x(50) & x(59) & x(73) & x(77) & x(80) & x(89) & x(102) & x(121) & x(136) & x(138) & x(142) & x(175) & x(177) & x(199) & x(221);
    y(11) <= not(p11_out);
    p11 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111100001000010000",
            TABLE => "0000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010011110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101101110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p11_in,
            y(0) => p11_out,
            y(1 to 14 - 1) => dummy11
        );


    p12_in <= x(3) & x(11) & x(22) & x(28) & x(29) & x(30) & x(42) & x(71) & x(113) & x(121) & x(162) & x(183) & x(202) & x(205) & x(236) & x(247) & x(253);
    y(12) <= not(p12_out);
    p12 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00100100110110101",
            TABLE => "11010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100101001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011001001101000001001101111101001101010011010010010011011011010011010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p12_in,
            y(0) => p12_out,
            y(1 to 14 - 1) => dummy12
        );


    p13_in <= x(16) & x(22) & x(26) & x(29) & x(43) & x(49) & x(54) & x(56) & x(58) & x(67) & x(76) & x(143) & x(204) & x(208) & x(217) & x(246);
    y(13) <= not(p13_out);
    p13 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110111011101011",
            TABLE => "0000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010001000001110001000110000111000110010110011010010000000000000000",
            SHIFT => 4,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p13_in,
            y(0) => p13_out,
            y(1 to 14 - 1) => dummy13
        );


    p14_in <= x(17) & x(18) & x(31) & x(51) & x(74) & x(99) & x(162) & x(171) & x(174) & x(183) & x(195);
    y(14) <= not(p14_out);
    p14 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01001001010",
            TABLE => "10110010001000001111101110110010001000000000000010110010001000001011001000100100110110111011001000100100010011011011001000100100100101100110100101101001100101100110100110010110100101100110100110110010111110110010000010110010101100101101101100100100101100101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p14_in,
            y(0) => p14_out,
            y(1 to 13 - 1) => dummy14
        );


    p15_in <= x(9) & x(14) & x(59) & x(84) & x(85) & x(114) & x(166) & x(238) & x(252) & x(253);
    y(15) <= not(p15_out);
    p15 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001101010",
            TABLE => "0010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100010000010110010001001001011001001101001100101100000000000000000",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p15_in,
            y(0) => p15_out,
            y(1 to 14 - 1) => dummy15
        );


    p16_in <= x(7) & x(18) & x(31) & x(38) & x(48) & x(66) & x(72) & x(85) & x(89) & x(98) & x(104) & x(106) & x(113) & x(133) & x(137) & x(154) & x(165) & x(173) & x(182) & x(209) & x(214) & x(220) & x(235) & x(239) & x(244) & x(251) & x(253);
    y(16) <= not(p16_out);
    p16 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011000110100001001001110111",
            TABLE => "100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p16_in,
            y(0) => p16_out,
            y(1 to 14 - 1) => dummy16
        );


    p17_in <= x(8) & x(23) & x(29) & x(31) & x(32) & x(53) & x(84) & x(95) & x(103) & x(107) & x(117) & x(118) & x(119) & x(125) & x(126) & x(132) & x(160) & x(181) & x(186) & x(201) & x(213) & x(228) & x(230) & x(244) & x(245);
    y(17) <= not(p17_out);
    p17 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110011111010111000110011",
            TABLE => "0100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p17_in,
            y(0) => p17_out,
            y(1 to 14 - 1) => dummy17
        );


    p18_in <= x(5) & x(6) & x(16) & x(27) & x(47) & x(51) & x(53) & x(68) & x(80) & x(100) & x(102) & x(103) & x(124) & x(132) & x(134) & x(140) & x(141) & x(147) & x(150) & x(177) & x(181) & x(186) & x(211) & x(240) & x(245);
    y(18) <= not(p18_out);
    p18 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111100001100000111011100",
            TABLE => "0000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p18_in,
            y(0) => p18_out,
            y(1 to 14 - 1) => dummy18
        );


    p19_in <= x(19) & x(28) & x(43) & x(50) & x(65) & x(88) & x(94) & x(97) & x(111) & x(119) & x(135) & x(158) & x(176) & x(189) & x(194) & x(199) & x(232) & x(252) & x(253) & x(255);
    y(19) <= not(p19_out);
    p19 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10111100000011010010",
            TABLE => "000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p19_in,
            y(0) => p19_out,
            y(1 to 14 - 1) => dummy19
        );


    p20_in <= x(38) & x(46) & x(48) & x(57) & x(60) & x(61) & x(63) & x(83) & x(105) & x(114) & x(117) & x(120) & x(123) & x(128) & x(154) & x(164) & x(189) & x(196) & x(216) & x(235) & x(238);
    y(20) <= not(p20_out);
    p20 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101010000111101100011",
            TABLE => "001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p20_in,
            y(0) => p20_out,
            y(1 to 14 - 1) => dummy20
        );


    p21_in <= x(11) & x(48) & x(107) & x(186) & x(213) & x(246);
    y(21) <= not(p21_out);
    p21 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101010",
            TABLE => "001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p21_in,
            y(0) => p21_out,
            y(1 to 13 - 1) => dummy21
        );


    p22_in <= x(5) & x(16) & x(19) & x(22) & x(47) & x(52) & x(63) & x(68) & x(80) & x(97) & x(110) & x(119) & x(120) & x(126) & x(142) & x(143) & x(164) & x(177) & x(181) & x(186) & x(223) & x(240) & x(251) & x(253);
    y(22) <= not(p22_out);
    p22 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001001011010110011001111",
            TABLE => "110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p22_in,
            y(0) => p22_out,
            y(1 to 14 - 1) => dummy22
        );


    p23_in <= x(11) & x(22) & x(28) & x(33) & x(57) & x(60) & x(63) & x(121) & x(138) & x(148) & x(152) & x(184) & x(189) & x(191) & x(194) & x(199) & x(208) & x(236) & x(248);
    y(23) <= not(p23_out);
    p23 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0101101111101001111",
            TABLE => "0010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101100000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p23_in,
            y(0) => p23_out,
            y(1 to 14 - 1) => dummy23
        );


    p24_in <= x(4) & x(48) & x(55) & x(57) & x(62) & x(77) & x(90) & x(99) & x(114) & x(144) & x(147) & x(176) & x(189) & x(194) & x(228) & x(241);
    y(24) <= not(p24_out);
    p24 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001000001011000",
            TABLE => "1110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101101101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010011000000011101000100000011110100010010110011010010000000000000000",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p24_in,
            y(0) => p24_out,
            y(1 to 14 - 1) => dummy24
        );


    p25_in <= x(0) & x(20) & x(186) & x(206) & x(241);
    y(25) <= not(p25_out);
    p25 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00010",
            TABLE => "11111011101100101011001000100000110110111011001010110010001001000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 5,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p25_in,
            y(0) => p25_out,
            y(1 to 13 - 1) => dummy25
        );


    p26_in <= x(14) & x(50) & x(57) & x(60) & x(61) & x(74) & x(91) & x(102) & x(106) & x(124) & x(140) & x(141) & x(148) & x(151) & x(155) & x(170) & x(172) & x(175) & x(202) & x(208) & x(229);
    y(26) <= not(p26_out);
    p26 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010101000110010010001",
            TABLE => "010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001110101001001011011111111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p26_in,
            y(0) => p26_out,
            y(1 to 14 - 1) => dummy26
        );


    p27_in <= x(14) & x(27) & x(44) & x(59) & x(85) & x(89) & x(125) & x(130) & x(175) & x(178) & x(179) & x(182) & x(194) & x(229) & x(253) & x(255);
    y(27) <= not(p27_out);
    p27 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110110101011001",
            TABLE => "0001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101100100000011010100010000101101010001101001100101100000000000000000",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p27_in,
            y(0) => p27_out,
            y(1 to 14 - 1) => dummy27
        );


    p28_in <= x(5) & x(28) & x(32) & x(47) & x(62) & x(65) & x(68) & x(70) & x(85) & x(102) & x(105) & x(106) & x(132) & x(140) & x(143) & x(146) & x(152) & x(177) & x(221) & x(232) & x(240) & x(248);
    y(28) <= not(p28_out);
    p28 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100101010001100011110",
            TABLE => "1011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010011000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101100000001000101011010000100010101110010110011010010000000000000000",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p28_in,
            y(0) => p28_out,
            y(1 to 14 - 1) => dummy28
        );


    p29_in <= x(2) & x(5) & x(6) & x(16) & x(37) & x(50) & x(67) & x(68) & x(70) & x(82) & x(84) & x(102) & x(113) & x(134) & x(151) & x(188) & x(189) & x(194) & x(247);
    y(29) <= not(p29_out);
    p29 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111000001010001011",
            TABLE => "0000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101101101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010011101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p29_in,
            y(0) => p29_out,
            y(1 to 14 - 1) => dummy29
        );


    p30_in <= x(19) & x(36) & x(50) & x(52) & x(82) & x(98) & x(125) & x(147) & x(160) & x(164) & x(165) & x(166) & x(168) & x(185) & x(208) & x(210) & x(211) & x(224) & x(229) & x(236) & x(238) & x(245) & x(246) & x(247);
    y(30) <= not(p30_out);
    p30 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000110110110101001110111",
            TABLE => "101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p30_in,
            y(0) => p30_out,
            y(1 to 14 - 1) => dummy30
        );


    p31_in <= x(15) & x(32) & x(46) & x(60) & x(62) & x(63) & x(89) & x(95) & x(154) & x(180) & x(216) & x(228) & x(235) & x(236) & x(238) & x(253) & x(255);
    y(31) <= not(p31_out);
    p31 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01100111001001001",
            TABLE => "01000000110101001101010011111101000000000100000001000000110101000100001011010100110101001011110100101011010000100100001011010100011010011001011010010110011010011001011001101001011010011001011000100000000000001011001000100000101100100010000011111011101100100010010001001101101100100010010010110010001001001101101110110010011010011001011010010110011010011001011001101001011010011001011011010100111111010100000011010100110101001011110101000010110101001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p31_in,
            y(0) => p31_out,
            y(1 to 14 - 1) => dummy31
        );


    p32_in <= x(35) & x(36) & x(40) & x(60) & x(76) & x(82) & x(112) & x(137) & x(138) & x(146) & x(153) & x(164) & x(165) & x(184) & x(187) & x(207) & x(235) & x(240) & x(244) & x(245);
    y(32) <= not(p32_out);
    p32 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10101110101110100111",
            TABLE => "000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p32_in,
            y(0) => p32_out,
            y(1 to 14 - 1) => dummy32
        );


    p33_in <= x(19) & x(44) & x(47) & x(51) & x(56) & x(58) & x(66) & x(71) & x(76) & x(91) & x(99) & x(107) & x(188) & x(195) & x(202) & x(213) & x(229) & x(247);
    y(33) <= not(p33_out);
    p33 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000110111010010011",
            TABLE => "101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p33_in,
            y(0) => p33_out,
            y(1 to 14 - 1) => dummy33
        );


    p34_in <= x(7) & x(30) & x(35) & x(40) & x(55) & x(60) & x(63) & x(65) & x(90) & x(102) & x(113) & x(117) & x(137) & x(139) & x(154) & x(161) & x(181) & x(184) & x(187) & x(196) & x(206) & x(207) & x(235) & x(253);
    y(34) <= not(p34_out);
    p34 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000001000000111001001110",
            TABLE => "111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p34_in,
            y(0) => p34_out,
            y(1 to 14 - 1) => dummy34
        );


    p35_in <= x(15) & x(19) & x(48) & x(55) & x(64) & x(72) & x(89) & x(111) & x(126) & x(179) & x(182) & x(189) & x(190) & x(193) & x(194) & x(216) & x(246) & x(252);
    y(35) <= not(p35_out);
    p35 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001100110010011111",
            TABLE => "100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p35_in,
            y(0) => p35_out,
            y(1 to 14 - 1) => dummy35
        );


    p36_in <= x(6) & x(8) & x(31) & x(54) & x(74) & x(77) & x(95) & x(117) & x(119) & x(121) & x(123) & x(131) & x(138) & x(190) & x(191) & x(198) & x(200) & x(202) & x(205) & x(232) & x(236) & x(238);
    y(36) <= not(p36_out);
    p36 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000111001011001010010",
            TABLE => "1111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101101011001000100000101100100010010010010110011010010000000000000000",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p36_in,
            y(0) => p36_out,
            y(1 to 14 - 1) => dummy36
        );


    p37_in <= x(1) & x(11) & x(14) & x(16) & x(24) & x(33) & x(38) & x(61) & x(63) & x(76) & x(77) & x(80) & x(123) & x(126) & x(142) & x(154) & x(158) & x(164) & x(166) & x(175) & x(183) & x(186) & x(188) & x(189) & x(196) & x(202) & x(238) & x(249) & x(253);
    y(37) <= not(p37_out);
    p37 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10011101110000101010010110010",
            TABLE => "00010111000000010000000100000000011111110001011100010111000000010001011110000001100000011110100001111110000101110001011110000001100101100110100101101001100101100110100110010110100101100110100100001000100011101000111011101111000000000000100000001000100011100001100010001110100011101110011101110001000110000001100010001110011010011001011010010110011010011001011001101001011010011001011010110010111110110010000010110010001000001011001000000000001000001011001011011011001001001011001000100100101100100100110100100100100101100110100101101001100101100110100110010110100101100110100101001101000001000000010000000000110111110100110101001101000001000100110100100100001001001011001011011011010011010100110100100100011010011001011010010110011010011001011001101001011010011001011010110010001000001111101110110010101100100010010011011011101100101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p37_in,
            y(0) => p37_out,
            y(1 to 14 - 1) => dummy37
        );


    p38_in <= x(11) & x(29) & x(55) & x(66) & x(71) & x(90) & x(91) & x(94) & x(96) & x(117) & x(158) & x(174) & x(179) & x(186) & x(195) & x(200) & x(213) & x(247);
    y(38) <= not(p38_out);
    p38 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110000101010000010",
            TABLE => "100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p38_in,
            y(0) => p38_out,
            y(1 to 14 - 1) => dummy38
        );


    p39_in <= x(8) & x(16) & x(53) & x(61) & x(77) & x(103) & x(109) & x(113) & x(115) & x(125) & x(126) & x(131) & x(138) & x(145) & x(148) & x(201) & x(217) & x(226) & x(242) & x(248);
    y(39) <= not(p39_out);
    p39 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101100011110010010",
            TABLE => "011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p39_in,
            y(0) => p39_out,
            y(1 to 14 - 1) => dummy39
        );


    p40_in <= x(55) & x(84) & x(87) & x(99) & x(108) & x(120) & x(128) & x(135) & x(178) & x(197) & x(223) & x(228) & x(234);
    y(40) <= not(p40_out);
    p40 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0101010001100",
            TABLE => "0100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101101011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p40_in,
            y(0) => p40_out,
            y(1 to 14 - 1) => dummy40
        );


    p41_in <= x(14) & x(17) & x(84) & x(91) & x(95) & x(112) & x(123) & x(161) & x(176) & x(201) & x(226) & x(228) & x(232) & x(236) & x(238);
    y(41) <= not(p41_out);
    p41 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100101100011101",
            TABLE => "010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110010011010110100111111111",
            SHIFT => 5,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p41_in,
            y(0) => p41_out,
            y(1 to 14 - 1) => dummy41
        );


    p42_in <= x(1) & x(6) & x(8) & x(17) & x(37) & x(39) & x(42) & x(51) & x(68) & x(94) & x(102) & x(103) & x(113) & x(117) & x(121) & x(132) & x(135) & x(140) & x(161) & x(167) & x(172) & x(182) & x(184) & x(187) & x(193) & x(219) & x(223) & x(225);
    y(42) <= not(p42_out);
    p42 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1011010110101110001011011111",
            TABLE => "0000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101100000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p42_in,
            y(0) => p42_out,
            y(1 to 14 - 1) => dummy42
        );


    p43_in <= x(1) & x(25) & x(28) & x(75) & x(78) & x(96) & x(101) & x(103) & x(107) & x(115) & x(118) & x(128) & x(174) & x(175) & x(190) & x(205) & x(211) & x(213) & x(223) & x(228) & x(238) & x(251);
    y(43) <= not(p43_out);
    p43 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111011110100000011001",
            TABLE => "0000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010011111110111010100110101000100000011010100010000000100000000000000101111011101010011010100010000101101010001000010010000100010101101101001100101101001011001101001100101100110100101101001100101100100000011010100010000101101010001101001100101100000000000000000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p43_in,
            y(0) => p43_out,
            y(1 to 14 - 1) => dummy43
        );


    p44_in <= x(5) & x(6) & x(40) & x(98) & x(121) & x(137) & x(138) & x(161) & x(164) & x(168) & x(185) & x(187) & x(235) & x(240) & x(244);
    y(44) <= not(p44_out);
    p44 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001010111101011",
            TABLE => "101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p44_in,
            y(0) => p44_out,
            y(1 to 13 - 1) => dummy44
        );


    p45_in <= x(14) & x(15) & x(16) & x(53) & x(59) & x(62) & x(72) & x(84) & x(89) & x(98) & x(115) & x(130) & x(138) & x(142) & x(171) & x(174) & x(175) & x(224);
    y(45) <= not(p45_out);
    p45 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110011100110100110",
            TABLE => "000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p45_in,
            y(0) => p45_out,
            y(1 to 14 - 1) => dummy45
        );


    p46_in <= x(3) & x(17) & x(20) & x(41) & x(64) & x(107) & x(109) & x(115) & x(119) & x(122) & x(124) & x(126) & x(133) & x(217) & x(231) & x(234) & x(237) & x(239);
    y(46) <= not(p46_out);
    p46 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100000111000001100",
            TABLE => "111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p46_in,
            y(0) => p46_out,
            y(1 to 14 - 1) => dummy46
        );


    p47_in <= x(5) & x(12) & x(47) & x(48) & x(55) & x(87) & x(88) & x(91) & x(93) & x(110) & x(112) & x(144) & x(151) & x(164) & x(172) & x(177) & x(188) & x(204) & x(206) & x(210) & x(255);
    y(47) <= not(p47_out);
    p47 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111001010011000010111",
            TABLE => "000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p47_in,
            y(0) => p47_out,
            y(1 to 14 - 1) => dummy47
        );


    p48_in <= x(7) & x(10) & x(42) & x(52) & x(55) & x(90) & x(94) & x(96) & x(105) & x(129) & x(139) & x(144) & x(147) & x(152) & x(153) & x(176) & x(178) & x(189) & x(207) & x(253) & x(254);
    y(48) <= not(p48_out);
    p48 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110111100100101010011",
            TABLE => "000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p48_in,
            y(0) => p48_out,
            y(1 to 14 - 1) => dummy48
        );


    p49_in <= x(8) & x(9) & x(19) & x(21) & x(38) & x(48) & x(55) & x(60) & x(74) & x(83) & x(120) & x(159) & x(164) & x(180) & x(182) & x(185) & x(190) & x(206) & x(210) & x(224) & x(233) & x(238) & x(245) & x(251);
    y(49) <= not(p49_out);
    p49 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000111101000101000011010",
            TABLE => "011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p49_in,
            y(0) => p49_out,
            y(1 to 14 - 1) => dummy49
        );


    p50_in <= x(26) & x(77) & x(97) & x(144) & x(178) & x(198) & x(229) & x(253) & x(255);
    y(50) <= not(p50_out);
    p50 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001110001",
            TABLE => "001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110110101001001011011111111",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p50_in,
            y(0) => p50_out,
            y(1 to 14 - 1) => dummy50
        );


    p51_in <= x(10) & x(36) & x(38) & x(53) & x(55) & x(61) & x(63) & x(83) & x(90) & x(106) & x(109) & x(110) & x(115) & x(117) & x(126) & x(144) & x(147) & x(155) & x(158) & x(160) & x(166) & x(185) & x(191) & x(197) & x(209) & x(216) & x(254);
    y(51) <= not(p51_out);
    p51 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111110001101011010000001101",
            TABLE => "000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110010011010110100111111111",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p51_in,
            y(0) => p51_out,
            y(1 to 14 - 1) => dummy51
        );


    p52_in <= x(3) & x(19) & x(21) & x(24) & x(38) & x(51) & x(65) & x(66) & x(98) & x(117) & x(122) & x(129) & x(131) & x(165) & x(168) & x(185) & x(193) & x(206) & x(208) & x(210) & x(217) & x(230) & x(231) & x(235) & x(239);
    y(52) <= not(p52_out);
    p52 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010111101101110101011001",
            TABLE => "0111000111110111000100000111000100010000011100010000000000010000011100011110011100011000011100010001100001110001100011100001100001101001100101101001011001101001100101100110100101101001100101100000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010010000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010010000100010001110000000000000100010001110111011110000100010001110000110001000111001110001000110001000111011100111000110001000111001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 3,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p52_in,
            y(0) => p52_out,
            y(1 to 13 - 1) => dummy52
        );


    p53_in <= x(18) & x(31) & x(48) & x(66) & x(67) & x(94) & x(96) & x(103) & x(132) & x(135) & x(149) & x(164) & x(176) & x(180) & x(214) & x(220) & x(221) & x(230) & x(239);
    y(53) <= not(p53_out);
    p53 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100101000101111100",
            TABLE => "0010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101101011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010010000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p53_in,
            y(0) => p53_out,
            y(1 to 14 - 1) => dummy53
        );


    p54_in <= x(0) & x(29) & x(98) & x(133) & x(137) & x(164) & x(165) & x(168) & x(182) & x(185) & x(193) & x(206) & x(208) & x(209) & x(217) & x(230) & x(235) & x(239) & x(247);
    y(54) <= not(p54_out);
    p54 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001011110101111011",
            TABLE => "0100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101100000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010010000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p54_in,
            y(0) => p54_out,
            y(1 to 14 - 1) => dummy54
        );


    p55_in <= x(5) & x(7) & x(23) & x(52) & x(55) & x(87) & x(90) & x(135) & x(158) & x(164) & x(176) & x(184) & x(189) & x(206) & x(220) & x(223) & x(232) & x(246) & x(251);
    y(55) <= not(p55_out);
    p55 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000010010101110000",
            TABLE => "1101010001000000010000000000000011111101110101001101010001000000110101000100001001000010001010111011110111010100110101000100001010010110011010010110100110010110011010011001011010010110011010011011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010010000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p55_in,
            y(0) => p55_out,
            y(1 to 14 - 1) => dummy55
        );


    p56_in <= x(14) & x(17) & x(42) & x(50) & x(112) & x(126) & x(134) & x(141) & x(151) & x(181) & x(189) & x(190) & x(194) & x(198) & x(201) & x(207) & x(226) & x(233) & x(234) & x(236) & x(241) & x(245) & x(255);
    y(56) <= not(p56_out);
    p56 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110110101001110101110",
            TABLE => "00000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100100100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011000000100010011010100110111011111000000000000010000000100010011010010010001001101010011011101101110110010001001000010010001001101100101100110100101101001100101100110100110010110100101100110100100101011101111110000001000101011001010111011110101000010001010110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p56_in,
            y(0) => p56_out,
            y(1 to 14 - 1) => dummy56
        );


    p57_in <= x(11) & x(16) & x(29) & x(36) & x(41);
    y(57) <= not(p57_out);
    p57 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01001",
            TABLE => "11010100111111010100000011010100110101001011110101000010110101001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 6,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p57_in,
            y(0) => p57_out,
            y(1 to 14 - 1) => dummy57
        );


    p58_in <= x(8) & x(16) & x(23) & x(33) & x(34) & x(41) & x(43) & x(51) & x(58) & x(116) & x(126) & x(132) & x(153) & x(202) & x(215) & x(249) & x(252);
    y(58) <= not(p58_out);
    p58 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11011011110000010",
            TABLE => "00000010000000000010101100000010001010110000001010111111001010110100001011010100001010110100001000101011010000101011110100101011100101100110100101101001100101100110100110010110100101100110100100000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100111111011101100101011001000100000110110111011001010110010001001000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p58_in,
            y(0) => p58_out,
            y(1 to 14 - 1) => dummy58
        );


    p59_in <= x(5) & x(8) & x(11) & x(16) & x(32) & x(35) & x(47) & x(65) & x(70) & x(88) & x(92) & x(132) & x(140) & x(141) & x(146) & x(164) & x(175) & x(180) & x(211) & x(223) & x(224) & x(232) & x(240);
    y(59) <= not(p59_out);
    p59 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00100100001110010001111",
            TABLE => "11010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100111110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100110001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100100010111011111110000000100010111000101110111111010000001000101111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p59_in,
            y(0) => p59_out,
            y(1 to 14 - 1) => dummy59
        );


    p60_in <= x(25) & x(39) & x(55) & x(69) & x(103) & x(107) & x(108) & x(113) & x(118) & x(119) & x(123) & x(149) & x(161) & x(162) & x(178) & x(181) & x(182) & x(193) & x(212) & x(234) & x(237) & x(250);
    y(60) <= not(p60_out);
    p60 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110001101011011111100",
            TABLE => "1000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100000100010001110000110001000111001101001100101100000000000000000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p60_in,
            y(0) => p60_out,
            y(1 to 14 - 1) => dummy60
        );


    p62_in <= x(0) & x(6) & x(16) & x(19) & x(36) & x(61) & x(77) & x(107) & x(190) & x(197) & x(206) & x(210) & x(212) & x(238);
    y(62) <= not(p62_out);
    p62 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000100000010",
            TABLE => "110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 5,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p62_in,
            y(0) => p62_out,
            y(1 to 14 - 1) => dummy62
        );


    p63_in <= x(24) & x(30) & x(40) & x(61) & x(66) & x(86) & x(94) & x(96) & x(97) & x(143) & x(154) & x(158) & x(164) & x(170) & x(177) & x(183) & x(184) & x(186) & x(213) & x(222) & x(227) & x(253);
    y(63) <= not(p63_out);
    p63 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001111011010100110010",
            TABLE => "0001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101101011001000100000101100100010010010010110011010010000000000000000",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p63_in,
            y(0) => p63_out,
            y(1 to 14 - 1) => dummy63
        );


    p64_in <= x(8) & x(22) & x(26) & x(30) & x(31) & x(38) & x(61) & x(74) & x(81) & x(83) & x(97) & x(99) & x(101) & x(115) & x(124) & x(131) & x(140) & x(160) & x(174) & x(211) & x(233) & x(237);
    y(64) <= not(p64_out);
    p64 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111010100001011100011",
            TABLE => "0000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010011110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010111000100010000011100010001100001101001100101100000000000000000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p64_in,
            y(0) => p64_out,
            y(1 to 14 - 1) => dummy64
        );


    p65_in <= x(8) & x(14) & x(22) & x(26) & x(32) & x(38) & x(47) & x(71) & x(74) & x(85) & x(91) & x(101) & x(110) & x(183) & x(208) & x(228);
    y(65) <= not(p65_out);
    p65 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000100100001010",
            TABLE => "1011001000100000001000000000000011111011101100101011001000100000101100100010010000100100010011011101101110110010101100100010010010010110011010010110100110010110011010011001011010010110011010011110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101100010000010110010001001001011001001101001100101100000000000000000",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p65_in,
            y(0) => p65_out,
            y(1 to 14 - 1) => dummy65
        );


    p66_in <= x(13) & x(14) & x(29) & x(42) & x(46) & x(73) & x(84) & x(94) & x(96) & x(114) & x(122) & x(123) & x(136) & x(149) & x(166) & x(180) & x(187) & x(207) & x(217) & x(247) & x(253);
    y(66) <= not(p66_out);
    p66 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101100101000011101000",
            TABLE => "000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001111010000110100111111111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p66_in,
            y(0) => p66_out,
            y(1 to 14 - 1) => dummy66
        );


    p67_in <= x(41) & x(197) & x(208) & x(234);
    y(67) <= not(p67_out);
    p67 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110",
            TABLE => "0000001000101011010000100010101110010110011010010000000000000000",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p67_in,
            y(0) => p67_out,
            y(1 to 14 - 1) => dummy67
        );


    p68_in <= x(1) & x(6) & x(9) & x(15) & x(19) & x(22) & x(25) & x(28) & x(33) & x(56) & x(60) & x(76) & x(104) & x(113) & x(122) & x(126) & x(131) & x(137) & x(139) & x(148) & x(171) & x(184) & x(193);
    y(68) <= not(p68_out);
    p68 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000100100111100001101",
            TABLE => "11010100010000000100000000000000111111011101010011010100010000001101010001000010010000100010101110111101110101001101010001000010100101100110100101101001100101100110100110010110100101100110100111010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100100000000100000001000000011101000100000001110100011101000111111100001011110000001100000011110100010000001111010001110100001111110011010011001011010010110011010011001011001101001011010011001011001001101110111110000010001001101010011011101101100100100010011010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p68_in,
            y(0) => p68_out,
            y(1 to 14 - 1) => dummy68
        );


    p69_in <= x(4) & x(25) & x(35) & x(44) & x(56) & x(57) & x(60) & x(89) & x(113) & x(126) & x(139) & x(148) & x(184) & x(196) & x(216) & x(255);
    y(69) <= not(p69_out);
    p69 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1011010110010111",
            TABLE => "0000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100001011100000001000101111000000110010110011010010000000000000000",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p69_in,
            y(0) => p69_out,
            y(1 to 14 - 1) => dummy69
        );


    p70_in <= x(8) & x(23) & x(31) & x(32) & x(38) & x(56) & x(73) & x(83) & x(97) & x(103) & x(106) & x(119) & x(125) & x(126) & x(132) & x(133) & x(160) & x(183) & x(191) & x(202) & x(249) & x(253);
    y(70) <= not(p70_out);
    p70 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100101001101111010101",
            TABLE => "1011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010010010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100100110100000100010011010010010001101001100101100000000000000000",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p70_in,
            y(0) => p70_out,
            y(1 to 14 - 1) => dummy70
        );


    p71_in <= x(5) & x(18) & x(29) & x(35) & x(37) & x(40) & x(45) & x(47) & x(50) & x(58) & x(62) & x(82) & x(83) & x(85) & x(112) & x(116) & x(121) & x(123) & x(133) & x(138) & x(139) & x(144) & x(153) & x(161) & x(164) & x(171) & x(179) & x(187) & x(212) & x(235) & x(238) & x(240) & x(244);
    y(71) <= not(p71_out);
    p71 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001101100011111110110011100110011",
            TABLE => "010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p71_in,
            y(0) => p71_out,
            y(1 to 15 - 1) => dummy71
        );


    p72_in <= x(1) & x(20) & x(33) & x(73) & x(74) & x(85) & x(103) & x(131) & x(144) & x(149) & x(163) & x(179) & x(192) & x(199) & x(208) & x(213) & x(215) & x(217) & x(224) & x(247) & x(250);
    y(72) <= not(p72_out);
    p72 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111100001001111001011",
            TABLE => "000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001011100010110100111111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p72_in,
            y(0) => p72_out,
            y(1 to 14 - 1) => dummy72
        );


    p73_in <= x(5) & x(8) & x(19) & x(47) & x(54) & x(75) & x(95) & x(103) & x(117) & x(119) & x(121) & x(123) & x(125) & x(126) & x(132) & x(133) & x(138) & x(141) & x(145) & x(178) & x(181) & x(194) & x(225) & x(228) & x(245);
    y(73) <= not(p73_out);
    p73 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010011100101111100000001",
            TABLE => "1101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010010010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101100000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p73_in,
            y(0) => p73_out,
            y(1 to 14 - 1) => dummy73
        );


    p74_in <= x(14) & x(20) & x(31) & x(37) & x(67) & x(73) & x(77) & x(80) & x(105) & x(106) & x(107) & x(112) & x(136) & x(138) & x(141) & x(167) & x(175) & x(192) & x(194) & x(202) & x(230) & x(231);
    y(74) <= not(p74_out);
    p74 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100011111111110101110",
            TABLE => "0100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010010000001000101011010000100010101110010110011010010000000000000000",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p74_in,
            y(0) => p74_out,
            y(1 to 14 - 1) => dummy74
        );


    p75_in <= x(8) & x(16) & x(31) & x(35) & x(41) & x(54) & x(58) & x(59) & x(73) & x(76) & x(89) & x(125) & x(126) & x(130) & x(138) & x(142) & x(191) & x(196) & x(202) & x(205) & x(249);
    y(75) <= not(p75_out);
    p75 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111101100110010111011",
            TABLE => "000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001011100010110100111111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p75_in,
            y(0) => p75_out,
            y(1 to 14 - 1) => dummy75
        );


    p76_in <= x(20) & x(77) & x(85) & x(125) & x(158) & x(163) & x(179) & x(189) & x(194) & x(207) & x(208) & x(210) & x(215) & x(238) & x(252);
    y(76) <= not(p76_out);
    p76 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011001001001111",
            TABLE => "010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 5,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p76_in,
            y(0) => p76_out,
            y(1 to 15 - 1) => dummy76
        );


    p77_in <= x(28) & x(31) & x(63) & x(65) & x(94) & x(96) & x(132) & x(135) & x(144) & x(145) & x(152) & x(172) & x(180) & x(194) & x(199) & x(204) & x(214) & x(216) & x(220) & x(255);
    y(77) <= not(p77_out);
    p77 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110100001110111010",
            TABLE => "000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p77_in,
            y(0) => p77_out,
            y(1 to 14 - 1) => dummy77
        );


    p78_in <= x(13) & x(14) & x(37) & x(50) & x(71) & x(73) & x(84) & x(122) & x(135) & x(136) & x(164) & x(166) & x(175) & x(198) & x(202) & x(217) & x(228) & x(248);
    y(78) <= not(p78_out);
    p78 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010001011110101111",
            TABLE => "110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p78_in,
            y(0) => p78_out,
            y(1 to 14 - 1) => dummy78
        );


    p79_in <= x(20) & x(55) & x(85) & x(98) & x(111) & x(120) & x(129) & x(131) & x(147) & x(179) & x(182) & x(189) & x(193) & x(202) & x(226) & x(246) & x(252);
    y(79) <= not(p79_out);
    p79 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01101001101011111",
            TABLE => "00100000101100101011001011111011000000000010000000100000101100100010010010110010101100101101101101001101001001000010010010110010011010011001011010010110011010011001011001101001011010011001011000100000101100101011001011111011000000000010000000100000101100100010010010110010101100101101101101001101001001000010010010110010011010011001011010010110011010011001011001101001011010011001011000000001000101110001011101111111100000010001011100010111011111100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p79_in,
            y(0) => p79_out,
            y(1 to 14 - 1) => dummy79
        );


    p80_in <= x(15) & x(34) & x(52) & x(69) & x(89) & x(125) & x(130) & x(135) & x(143) & x(152) & x(173) & x(176) & x(247) & x(251);
    y(80) <= not(p80_out);
    p80 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10110101001011",
            TABLE => "000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p80_in,
            y(0) => p80_out,
            y(1 to 13 - 1) => dummy80
        );


    p81_in <= x(14) & x(17) & x(24) & x(33) & x(59) & x(63) & x(71) & x(73) & x(80) & x(91) & x(103) & x(107) & x(112) & x(133) & x(138) & x(142) & x(159) & x(186) & x(188) & x(202) & x(207);
    y(81) <= not(p81_out);
    p81 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001101100000000101001",
            TABLE => "010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001110101001001011011111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p81_in,
            y(0) => p81_out,
            y(1 to 14 - 1) => dummy81
        );


    p82_in <= x(10) & x(17) & x(18) & x(20) & x(37) & x(41) & x(126) & x(163) & x(169) & x(181) & x(184) & x(191) & x(196) & x(225) & x(230) & x(236) & x(255);
    y(82) <= not(p82_out);
    p82 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11011110101000110",
            TABLE => "00000001000000000001011100000001000101110000000101111111000101111000000111101000000101111000000100010111100000010111111000010111011010011001011010010110011010011001011001101001011010011001011000100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011010111111001010110010101100000010101111010010101100101011010000101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p82_in,
            y(0) => p82_out,
            y(1 to 14 - 1) => dummy82
        );


    p83_in <= x(11) & x(20) & x(28) & x(33) & x(35) & x(46) & x(51) & x(62) & x(65) & x(66) & x(88) & x(96) & x(113) & x(122) & x(133) & x(137) & x(150) & x(163) & x(165) & x(186) & x(204) & x(210);
    y(83) <= not(p83_out);
    p83 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010000100010001110001",
            TABLE => "1000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010011101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010010111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101101101010001000000110101000100001010010110011010010000000000000000",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p83_in,
            y(0) => p83_out,
            y(1 to 14 - 1) => dummy83
        );


    p84_in <= x(3) & x(6) & x(28) & x(39) & x(42) & x(55) & x(62) & x(68) & x(80) & x(94) & x(96) & x(113) & x(121) & x(133) & x(135) & x(145) & x(158) & x(161) & x(172) & x(177) & x(193) & x(202) & x(206) & x(219) & x(230) & x(247) & x(250) & x(253);
    y(84) <= not(p84_out);
    p84 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001010110111100011111011001",
            TABLE => "1101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010010001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101100000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100100000011010100010000101101010001101001100101100000000000000000",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p84_in,
            y(0) => p84_out,
            y(1 to 14 - 1) => dummy84
        );


    p85_in <= x(41) & x(49) & x(54) & x(80) & x(84) & x(105) & x(119) & x(138) & x(191) & x(194) & x(201) & x(202) & x(232) & x(236) & x(238) & x(255);
    y(85) <= not(p85_out);
    p85 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001110100110100",
            TABLE => "0001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101101000111000001000100011100001100010010110011010010000000000000000",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p85_in,
            y(0) => p85_out,
            y(1 to 14 - 1) => dummy85
        );


    p86_in <= x(21) & x(24) & x(46) & x(59) & x(68) & x(73) & x(75) & x(87) & x(88) & x(94) & x(115) & x(117) & x(132) & x(140) & x(152) & x(167) & x(176) & x(178) & x(180) & x(186) & x(196) & x(226) & x(234) & x(237) & x(238) & x(254);
    y(86) <= not(p86_out);
    p86 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11100001010011010101110101",
            TABLE => "000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p86_in,
            y(0) => p86_out,
            y(1 to 14 - 1) => dummy86
        );


    p87_in <= x(4) & x(11) & x(26) & x(35) & x(38) & x(40) & x(45) & x(47) & x(51) & x(70) & x(74) & x(80) & x(81) & x(82) & x(83) & x(86) & x(100) & x(110) & x(132) & x(140) & x(146) & x(149) & x(152) & x(196) & x(202) & x(203) & x(221) & x(240) & x(244);
    y(87) <= not(p87_out);
    p87 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11010110100111100111000100111",
            TABLE => "00000100000000000100110100000100010011010000010011011111010011010010010010110010010011010010010001001101001001001101101101001101100101100110100101101001100101100110100110010110100101100110100101000000110101000000000001000000110101001111110101000000110101000100001011010100001010110100001011010100101111010100001011010100011010011001011010010110011010011001011001101001011010011001011000000000010000000100000011010100010000001101010011010100111111010010101101000010010000101101010001000010110101001101010010111101100101100110100101101001100101100110100110010110100101100110100101000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011001111111000101110001011100000001011111100001011100010111100000010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p87_in,
            y(0) => p87_out,
            y(1 to 14 - 1) => dummy87
        );


    p88_in <= x(8) & x(14) & x(16) & x(24) & x(32) & x(48) & x(78) & x(87) & x(97) & x(117) & x(123) & x(144) & x(147) & x(152) & x(200) & x(204) & x(208) & x(211) & x(213);
    y(88) <= not(p88_out);
    p88 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100000100010100101",
            TABLE => "1110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101101101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010011011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p88_in,
            y(0) => p88_out,
            y(1 to 14 - 1) => dummy88
        );


    p89_in <= x(11) & x(43) & x(48) & x(52) & x(55) & x(57) & x(61) & x(65) & x(72) & x(74) & x(85) & x(90) & x(91) & x(99) & x(120) & x(125) & x(134) & x(138) & x(144) & x(147) & x(153) & x(164) & x(168) & x(172) & x(182) & x(190) & x(210) & x(213) & x(224) & x(229) & x(233) & x(236) & x(238) & x(244) & x(245);
    y(89) <= not(p89_out);
    p89 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11000110101010101010000001110000100",
            TABLE => "01000000000000001101010001000000110101000100000011111101110101000100001000101011110101000100001011010100010000101011110111010100011010011001011010010110011010011001011001101001011010011001011000100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011000100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011011101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011000001000100011101000111011101111000000000000100000001000100011100001100010001110100011101110011101110001000110000001100010001110011010011001011010010110011010011001011001101001011010011001011011101111100011101000111000001000111001111000111010001110000110000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p89_in,
            y(0) => p89_out,
            y(1 to 14 - 1) => dummy89
        );


    p90_in <= x(58) & x(87) & x(99) & x(160) & x(178) & x(223);
    y(90) <= not(p90_out);
    p90 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001101",
            TABLE => "010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p90_in,
            y(0) => p90_out,
            y(1 to 13 - 1) => dummy90
        );


    p91_in <= x(33) & x(57) & x(60) & x(61) & x(63) & x(117) & x(123) & x(139) & x(154) & x(180) & x(196) & x(216) & x(235) & x(238);
    y(91) <= not(p91_out);
    p91 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11011000001100",
            TABLE => "000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p91_in,
            y(0) => p91_out,
            y(1 to 13 - 1) => dummy91
        );


    p92_in <= x(17) & x(18) & x(26) & x(29) & x(38) & x(47) & x(56) & x(58) & x(74) & x(99) & x(123) & x(158) & x(171);
    y(92) <= not(p92_out);
    p92 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001001001010",
            TABLE => "1000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010010100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p92_in,
            y(0) => p92_out,
            y(1 to 13 - 1) => dummy92
        );


    p93_in <= x(14) & x(30) & x(36) & x(78) & x(84) & x(106) & x(118) & x(119) & x(120) & x(122) & x(131) & x(132) & x(133) & x(137) & x(140) & x(150) & x(165) & x(183) & x(197) & x(222) & x(234) & x(237) & x(245);
    y(93) <= not(p93_out);
    p93 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11001110110110101111011",
            TABLE => "00010000000000000111000100010000011100010001000011110111011100010001100010001110011100010001100001110001000110001110011101110001100101100110100101101001100101100110100110010110100101100110100100000100010011010000000000000100010011011101111100000100010011010010010001001101101100100010010001001101110110110010010001001101100101100110100101101001100101100110100110010110100101100110100100010000011100010000000000010000011100011111011100010000011100010001100001110001100011100001100001110001111001110001100001110001100101100110100101101001100101100110100110010110100101100110100100010000011100010111000111110111000110000111000101110001111001111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p93_in,
            y(0) => p93_out,
            y(1 to 14 - 1) => dummy93
        );


    p94_in <= x(7) & x(12) & x(30) & x(33) & x(36) & x(60) & x(63) & x(88) & x(93) & x(107) & x(122) & x(168) & x(171) & x(184) & x(189) & x(190) & x(196) & x(204) & x(215) & x(233) & x(236);
    y(94) <= not(p94_out);
    p94 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010011000100010100100",
            TABLE => "011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001100011101001011011111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p94_in,
            y(0) => p94_out,
            y(1 to 14 - 1) => dummy94
        );


    p95_in <= x(15) & x(23) & x(60) & x(89) & x(115) & x(140) & x(175) & x(180) & x(211) & x(216) & x(232) & x(238) & x(245) & x(255);
    y(95) <= not(p95_out);
    p95 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10101011100100",
            TABLE => "001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p95_in,
            y(0) => p95_out,
            y(1 to 14 - 1) => dummy95
        );


    p96_in <= x(15) & x(20) & x(38) & x(48) & x(53) & x(72) & x(74) & x(80) & x(88) & x(111) & x(130) & x(171) & x(174) & x(180) & x(185) & x(220) & x(224) & x(232) & x(233) & x(252);
    y(96) <= not(p96_out);
    p96 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00111010011100001111",
            TABLE => "001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p96_in,
            y(0) => p96_out,
            y(1 to 14 - 1) => dummy96
        );


    p97_in <= x(14) & x(18) & x(43) & x(56) & x(71) & x(72) & x(91) & x(92) & x(111) & x(123) & x(134) & x(136) & x(143) & x(147) & x(151) & x(192) & x(194) & x(207) & x(213) & x(241);
    y(97) <= not(p97_out);
    p97 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11100110011100000110",
            TABLE => "000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p97_in,
            y(0) => p97_out,
            y(1 to 14 - 1) => dummy97
        );


    p98_in <= x(15) & x(48) & x(181) & x(186);
    y(98) <= not(p98_out);
    p98 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111",
            TABLE => "0001011100000001000101111000000110010110011010010000000000000000",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p98_in,
            y(0) => p98_out,
            y(1 to 13 - 1) => dummy98
        );


    p99_in <= x(11) & x(26) & x(88) & x(93) & x(94) & x(107) & x(112) & x(117) & x(132) & x(152) & x(172) & x(176) & x(181) & x(198) & x(226) & x(232) & x(237) & x(255);
    y(99) <= not(p99_out);
    p99 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100011101000001111",
            TABLE => "011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p99_in,
            y(0) => p99_out,
            y(1 to 14 - 1) => dummy99
        );


    p100_in <= x(5) & x(11) & x(16) & x(22) & x(23) & x(28) & x(50) & x(65) & x(88) & x(112) & x(179) & x(197) & x(203) & x(240) & x(252) & x(255);
    y(100) <= not(p100_out);
    p100 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100110001000111",
            TABLE => "0111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101101110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100001011100000001000101111000000110010110011010010000000000000000",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p100_in,
            y(0) => p100_out,
            y(1 to 14 - 1) => dummy100
        );


    p101_in <= x(16) & x(18) & x(19) & x(23) & x(33) & x(41) & x(58) & x(59) & x(60) & x(63) & x(76) & x(89) & x(125) & x(126) & x(142) & x(145) & x(147) & x(180) & x(202) & x(215) & x(249);
    y(101) <= not(p101_out);
    p101 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001101011000110011110",
            TABLE => "010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001001010110110100111111111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p101_in,
            y(0) => p101_out,
            y(1 to 14 - 1) => dummy101
        );


    p102_in <= x(17) & x(40) & x(50) & x(58) & x(70) & x(74) & x(80) & x(82) & x(83) & x(91) & x(99) & x(112) & x(123) & x(138) & x(139) & x(187) & x(192) & x(233) & x(244);
    y(102) <= not(p102_out);
    p102 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100001111110101001",
            TABLE => "1000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010010000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011000111000001000111011111000111000001000000000001000111000001000100011100001100011100111100011100001100001110001100011100001100010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p102_in,
            y(0) => p102_out,
            y(1 to 14 - 1) => dummy102
        );


    p103_in <= x(8) & x(31) & x(41) & x(69) & x(77) & x(165) & x(185) & x(197) & x(208);
    y(103) <= not(p103_out);
    p103 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110000100",
            TABLE => "100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001100011101001011011111111",
            SHIFT => 5,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p103_in,
            y(0) => p103_out,
            y(1 to 14 - 1) => dummy103
        );


    p104_in <= x(13) & x(14) & x(18) & x(19) & x(24) & x(41) & x(44) & x(71) & x(82) & x(84) & x(90) & x(91) & x(92) & x(99) & x(110) & x(112) & x(123) & x(125) & x(126) & x(135) & x(145) & x(154) & x(155) & x(176) & x(213) & x(219) & x(223) & x(245);
    y(104) <= not(p104_out);
    p104 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110001010010001100111101000",
            TABLE => "1000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101101011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010010000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010011000000011101000100000011110100010010110011010010000000000000000",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p104_in,
            y(0) => p104_out,
            y(1 to 14 - 1) => dummy104
        );


    p105_in <= x(14) & x(112) & x(135) & x(152) & x(163) & x(166) & x(176) & x(180) & x(186) & x(206) & x(228) & x(247);
    y(105) <= not(p105_out);
    p105 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000111110100",
            TABLE => "011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p105_in,
            y(0) => p105_out,
            y(1 to 13 - 1) => dummy105
        );


    p106_in <= x(8) & x(14) & x(23) & x(27) & x(29) & x(31) & x(43) & x(49) & x(50) & x(53) & x(61) & x(65) & x(70) & x(88) & x(89) & x(95) & x(103) & x(104) & x(112) & x(121) & x(132) & x(142) & x(164) & x(180) & x(194) & x(207) & x(232) & x(244);
    y(106) <= not(p106_out);
    p106 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110100001000011111110101011",
            TABLE => "0010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101101110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010000000000100000001000001011001000100000101100101011001011111011010011010010010000100100101100100010010010110010101100101101101110010110011010010110100110010110011010011001011010010110011010010001000001110001000110000111000110010110011010010000000000000000",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p106_in,
            y(0) => p106_out,
            y(1 to 14 - 1) => dummy106
        );


    p107_in <= x(3) & x(17) & x(20) & x(24) & x(41) & x(62) & x(69) & x(70) & x(113) & x(122) & x(137) & x(163) & x(208) & x(214) & x(217) & x(230) & x(231) & x(248);
    y(107) <= not(p107_out);
    p107 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100101000011010010",
            TABLE => "010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p107_in,
            y(0) => p107_out,
            y(1 to 14 - 1) => dummy107
        );


    p108_in <= x(3) & x(4) & x(26) & x(45) & x(60) & x(97) & x(112) & x(125) & x(172) & x(176) & x(203) & x(226) & x(253) & x(255);
    y(108) <= not(p108_out);
    p108 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11010110000101",
            TABLE => "000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p108_in,
            y(0) => p108_out,
            y(1 to 13 - 1) => dummy108
        );


    p109_in <= x(13) & x(49) & x(53) & x(60) & x(71) & x(75) & x(84) & x(95) & x(115) & x(171) & x(190) & x(197) & x(208) & x(217) & x(218) & x(228) & x(234) & x(237) & x(238) & x(241) & x(242) & x(246);
    y(109) <= not(p109_out);
    p109 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010111101011010010110",
            TABLE => "0001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010010000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p109_in,
            y(0) => p109_out,
            y(1 to 14 - 1) => dummy109
        );


    p110_in <= x(13) & x(14) & x(20) & x(32) & x(54) & x(71) & x(82) & x(84) & x(87) & x(88) & x(110) & x(112) & x(119) & x(126) & x(134) & x(157) & x(164) & x(174) & x(189) & x(190) & x(194) & x(195) & x(228) & x(232) & x(241) & x(246);
    y(110) <= not(p110_out);
    p110 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10110101011001110110010010",
            TABLE => "000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p110_in,
            y(0) => p110_out,
            y(1 to 14 - 1) => dummy110
        );


    p111_in <= x(2) & x(8) & x(11) & x(22) & x(31) & x(33) & x(36) & x(74) & x(78) & x(125) & x(132) & x(144) & x(159) & x(160) & x(171) & x(183) & x(194) & x(197) & x(199) & x(207) & x(225) & x(236) & x(248);
    y(111) <= not(p111_out);
    p111 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10010101011000110111011",
            TABLE => "01001101000001000000010000000000110111110100110101001101000001000100110100100100001001001011001011011011010011010100110100100100011010011001011010010110011010011001011001101001011010011001011000101011000000101011111100101011000000100000000000101011000000100010101101000010101111010010101101000010110101000010101101000010011010011001011010010110011010011001011001101001011010011001011001001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011000010000011100010111000111110111000110000111000101110001111001111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p111_in,
            y(0) => p111_out,
            y(1 to 14 - 1) => dummy111
        );


    p112_in <= x(8) & x(10) & x(18) & x(58) & x(61) & x(69) & x(77) & x(101) & x(116) & x(126) & x(131) & x(142) & x(144) & x(147) & x(170) & x(202) & x(213) & x(214) & x(241);
    y(112) <= not(p112_out);
    p112 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100011001100111001",
            TABLE => "1101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010010010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100000100010001110100011101110111100000000000010000000100010001110000110001000111010001110111001110111000100011000000110001000111001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p112_in,
            y(0) => p112_out,
            y(1 to 14 - 1) => dummy112
        );


    p113_in <= x(1) & x(13) & x(14) & x(25) & x(45) & x(56) & x(75) & x(76) & x(83) & x(96) & x(97) & x(101) & x(107) & x(108) & x(111) & x(115) & x(123) & x(126) & x(142) & x(146) & x(153) & x(194) & x(201) & x(234);
    y(113) <= not(p113_out);
    p113 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101011011010011100001101",
            TABLE => "000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p113_in,
            y(0) => p113_out,
            y(1 to 14 - 1) => dummy113
        );


    p114_in <= x(6) & x(17) & x(27) & x(35) & x(40) & x(51) & x(84) & x(89) & x(100) & x(119) & x(122) & x(124) & x(131) & x(133) & x(137) & x(138) & x(150) & x(165) & x(177) & x(178) & x(181) & x(228) & x(231) & x(234) & x(237) & x(240);
    y(114) <= not(p114_out);
    p114 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01011111001101010110000011",
            TABLE => "000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110111010001000000010000000000000001111111011101000111010001000000011101000100000011000000100010111011111101110100011101000100000010110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p114_in,
            y(0) => p114_out,
            y(1 to 14 - 1) => dummy114
        );


    p115_in <= x(14) & x(18) & x(21) & x(46) & x(59) & x(61) & x(84) & x(89) & x(103) & x(105) & x(107) & x(127) & x(132) & x(173) & x(175) & x(177) & x(186) & x(191) & x(197) & x(221) & x(222) & x(234) & x(235) & x(237) & x(250) & x(251);
    y(115) <= not(p115_out);
    p115 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00110011111010001010000110",
            TABLE => "100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p115_in,
            y(0) => p115_out,
            y(1 to 14 - 1) => dummy115
        );


    p116_in <= x(36) & x(54) & x(56) & x(75) & x(93) & x(95) & x(138) & x(228);
    y(116) <= not(p116_out);
    p116 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11001001",
            TABLE => "001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p116_in,
            y(0) => p116_out,
            y(1 to 13 - 1) => dummy116
        );


    p117_in <= x(0) & x(19) & x(25) & x(60) & x(63) & x(76) & x(113) & x(126) & x(148) & x(158) & x(176) & x(180) & x(181) & x(184) & x(193) & x(206) & x(212) & x(226) & x(235);
    y(117) <= not(p117_out);
    p117 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000111011001010110",
            TABLE => "0111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101100000100010001110000000000000100010001110111011110000100010001110000110001000111001110001000110001000111011100111000110001000111001101001100101101001011001101001100101100110100101101001100101100001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p117_in,
            y(0) => p117_out,
            y(1 to 14 - 1) => dummy117
        );


    p118_in <= x(27) & x(41) & x(63) & x(66) & x(77) & x(85) & x(135) & x(149) & x(212) & x(214) & x(230) & x(231) & x(239);
    y(118) <= not(p118_out);
    p118 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010010111010",
            TABLE => "0100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 5,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p118_in,
            y(0) => p118_out,
            y(1 to 14 - 1) => dummy118
        );


    p119_in <= x(11) & x(22) & x(43) & x(79) & x(80) & x(83) & x(88) & x(93) & x(112) & x(134) & x(135) & x(166) & x(172) & x(177) & x(179) & x(182) & x(236) & x(253) & x(254);
    y(119) <= not(p119_out);
    p119 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110101101101110111",
            TABLE => "0010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101100000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010010000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p119_in,
            y(0) => p119_out,
            y(1 to 14 - 1) => dummy119
        );


    p120_in <= x(6) & x(14) & x(20) & x(33) & x(35) & x(38) & x(40) & x(55) & x(72) & x(74) & x(80) & x(111) & x(120) & x(129) & x(131) & x(150) & x(154) & x(187) & x(194) & x(196) & x(224) & x(246) & x(251);
    y(120) <= not(p120_out);
    p120 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000101010100111010110",
            TABLE => "11010100010000000100000000000000111111011101010011010100010000001101010001000010010000100010101110111101110101001101010001000010100101100110100101101001100101100110100110010110100101100110100101001101000001001101111101001101000001000000000001001101000001000100110100100100110110110100110100100100101100100100110100100100011010011001011010010110011010011001011001101001011010011001011000101011101111110000001000101011000000100010101100000000000000100010101110111101010000100010101101000010001010111101010001000010011010011001011010010110011010011001011001101001011010011001011000101011000000101011111100101011001010110100001010111101001010110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p120_in,
            y(0) => p120_out,
            y(1 to 14 - 1) => dummy120
        );


    p121_in <= x(17) & x(28) & x(32) & x(51) & x(65) & x(74) & x(87) & x(117) & x(140) & x(162) & x(171) & x(185) & x(189) & x(214) & x(253);
    y(121) <= not(p121_out);
    p121 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010001101010100",
            TABLE => "110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110100011101001011011111111",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p121_in,
            y(0) => p121_out,
            y(1 to 13 - 1) => dummy121
        );


    p122_in <= x(5) & x(6) & x(9) & x(24) & x(40) & x(51) & x(56) & x(58) & x(61) & x(68) & x(80) & x(106) & x(126) & x(142) & x(177) & x(186) & x(187) & x(202) & x(203) & x(240) & x(244) & x(254);
    y(122) <= not(p122_out);
    p122 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000111001101010110110",
            TABLE => "1111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010010010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p122_in,
            y(0) => p122_out,
            y(1 to 14 - 1) => dummy122
        );


    p123_in <= x(17) & x(18) & x(62) & x(74) & x(126) & x(153) & x(162) & x(173) & x(177) & x(212) & x(230) & x(239);
    y(123) <= not(p123_out);
    p123 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011101011100",
            TABLE => "000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p123_in,
            y(0) => p123_out,
            y(1 to 14 - 1) => dummy123
        );


    p124_in <= x(4) & x(26) & x(46) & x(52) & x(60) & x(94) & x(96) & x(116) & x(125) & x(132) & x(140) & x(152) & x(176) & x(177) & x(186) & x(197) & x(223) & x(225) & x(226) & x(237) & x(251) & x(254);
    y(124) <= not(p124_out);
    p124 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010010101100011001101",
            TABLE => "0100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101101000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010000010001001101001001000100110110010110011010010000000000000000",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p124_in,
            y(0) => p124_out,
            y(1 to 14 - 1) => dummy124
        );


    p125_in <= x(19) & x(50) & x(55) & x(84) & x(111) & x(112) & x(129) & x(135) & x(158) & x(164) & x(168) & x(176) & x(178) & x(180) & x(182) & x(189) & x(193) & x(194) & x(198) & x(203) & x(220) & x(232) & x(239);
    y(125) <= not(p125_out);
    p125 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101101011010101100011",
            TABLE => "01110001111101110001000001110001000100000111000100000000000100000111000111100111000110000111000100011000011100011000111000011000011010011001011010010110011010011001011001101001011010011001011000101011000000101011111100101011000000100000000000101011000000100010101101000010101111010010101101000010110101000010101101000010011010011001011010010110011010011001011001101001011010011001011000010000011100010000000000010000011100011111011100010000011100010001100001110001100011100001100001110001111001110001100001110001100101100110100101101001100101100110100110010110100101100110100111110111011100010111000100010000111001110111000101110001000110001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p125_in,
            y(0) => p125_out,
            y(1 to 14 - 1) => dummy125
        );


    p126_in <= x(1) & x(25) & x(28) & x(33) & x(37) & x(45) & x(47) & x(52) & x(62) & x(65) & x(68) & x(70) & x(89) & x(100) & x(113) & x(120) & x(128) & x(146) & x(153) & x(173) & x(181) & x(199) & x(213) & x(221) & x(230) & x(239) & x(254);
    y(126) <= not(p126_out);
    p126 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100100100101111011001100111",
            TABLE => "100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 4,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p126_in,
            y(0) => p126_out,
            y(1 to 14 - 1) => dummy126
        );


    p127_in <= x(6) & x(29) & x(38) & x(40) & x(49) & x(50) & x(60) & x(83) & x(107) & x(108) & x(109) & x(120) & x(123) & x(133) & x(139) & x(153) & x(161) & x(187) & x(200) & x(212) & x(215) & x(221) & x(233) & x(234) & x(235);
    y(127) <= not(p127_out);
    p127 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0101000101100101110101010",
            TABLE => "1000111000001000111011111000111000001000000000001000111000001000100011100001100011100111100011100001100001110001100011100001100010010110011010010110100110010110011010011001011010010110011010010010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101100001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010010100110100000100110111110100110100000100000000000100110100000100010011010010010011011011010011010010010010110010010011010010010001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p127_in,
            y(0) => p127_out,
            y(1 to 14 - 1) => dummy127
        );


    p128_in <= x(13) & x(21) & x(25) & x(31) & x(38) & x(41) & x(55) & x(72) & x(83) & x(98) & x(106) & x(111) & x(122) & x(129) & x(131) & x(154) & x(160) & x(165) & x(166) & x(202) & x(209) & x(210) & x(217) & x(228) & x(236);
    y(128) <= not(p128_out);
    p128 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100111000111011010110111",
            TABLE => "0111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101100111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101100000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p128_in,
            y(0) => p128_out,
            y(1 to 14 - 1) => dummy128
        );


    p129_in <= x(3) & x(11) & x(24) & x(29) & x(38) & x(56) & x(58) & x(62) & x(99) & x(113) & x(122) & x(123) & x(141) & x(144) & x(145) & x(146) & x(147) & x(153) & x(244) & x(248);
    y(129) <= not(p129_out);
    p129 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001010011111110001",
            TABLE => "111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p129_in,
            y(0) => p129_out,
            y(1 to 14 - 1) => dummy129
        );


    p130_in <= x(0) & x(15) & x(19) & x(25) & x(46) & x(60) & x(64) & x(120) & x(123) & x(126) & x(128) & x(180) & x(186) & x(208) & x(226) & x(238) & x(241);
    y(130) <= not(p130_out);
    p130 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10001000001011101",
            TABLE => "10110010001000000010000000000000111110111011001010110010001000001011001000100100001001000100110111011011101100101011001000100100100101100110100101101001100101100110100110010110100101100110100111111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011000000100010011010100110111011111001001000100110101001101110110111001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p130_in,
            y(0) => p130_out,
            y(1 to 14 - 1) => dummy130
        );


    p131_in <= x(1) & x(3) & x(25) & x(78) & x(84) & x(92) & x(103) & x(107) & x(108) & x(115) & x(118) & x(120) & x(123) & x(128) & x(132) & x(134) & x(143) & x(178) & x(181) & x(194) & x(205) & x(211) & x(213) & x(223) & x(228) & x(234) & x(239) & x(251);
    y(131) <= not(p131_out);
    p131 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101010011000100111111001110",
            TABLE => "0000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010011000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101100000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010000001000101011010000100010101110010110011010010000000000000000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p131_in,
            y(0) => p131_out,
            y(1 to 14 - 1) => dummy131
        );


    p132_in <= x(0) & x(4) & x(35) & x(60) & x(64) & x(76) & x(82) & x(122) & x(132) & x(137) & x(146) & x(150) & x(164) & x(176) & x(180) & x(213) & x(235) & x(238) & x(247) & x(254);
    y(132) <= not(p132_out);
    p132 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11100111100010010011",
            TABLE => "000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p132_in,
            y(0) => p132_out,
            y(1 to 14 - 1) => dummy132
        );


    p133_in <= x(26) & x(30) & x(38) & x(70) & x(74) & x(116) & x(119) & x(121) & x(138) & x(152) & x(158) & x(162) & x(171) & x(183) & x(191) & x(197) & x(199) & x(203) & x(232) & x(233) & x(247);
    y(133) <= not(p133_out);
    p133 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111110011110110111010",
            TABLE => "000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p133_in,
            y(0) => p133_out,
            y(1 to 14 - 1) => dummy133
        );


    p134_in <= x(96) & x(152) & x(168) & x(185) & x(203) & x(206) & x(247);
    y(134) <= not(p134_out);
    p134 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0010001",
            TABLE => "1110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 5,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p134_in,
            y(0) => p134_out,
            y(1 to 13 - 1) => dummy134
        );


    p135_in <= x(0) & x(4) & x(6) & x(14) & x(20) & x(33) & x(35) & x(36) & x(38) & x(60) & x(69) & x(79) & x(81) & x(111) & x(129) & x(154) & x(173) & x(184) & x(196) & x(236) & x(247) & x(251) & x(253);
    y(135) <= not(p135_out);
    p135 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11011110001010101011111",
            TABLE => "00000001000000000001011100000001000101110000000101111111000101111000000111101000000101111000000100010111100000010111111000010111011010011001011010010110011010011001011001101001011010011001011010110010001000000010000000000000111110111011001010110010001000001011001000100100001001000100110111011011101100101011001000100100100101100110100101101001100101100110100110010110100101100110100100100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011000000001000101110001011101111111100000010001011100010111011111100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p135_in,
            y(0) => p135_out,
            y(1 to 14 - 1) => dummy135
        );


    p136_in <= x(24) & x(37) & x(38) & x(45) & x(50) & x(53) & x(70) & x(98) & x(102) & x(103) & x(118) & x(130) & x(138) & x(139) & x(170) & x(171) & x(185) & x(195) & x(203) & x(207) & x(247);
    y(136) <= not(p136_out);
    p136 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100100011000101011001",
            TABLE => "100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001110101001001011011111111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p136_in,
            y(0) => p136_out,
            y(1 to 14 - 1) => dummy136
        );


    p137_in <= x(8) & x(36) & x(61) & x(121) & x(133) & x(138) & x(191) & x(208) & x(241) & x(245);
    y(137) <= not(p137_out);
    p137 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001110111",
            TABLE => "0111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100001011100000001000101111000000110010110011010010000000000000000",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p137_in,
            y(0) => p137_out,
            y(1 to 14 - 1) => dummy137
        );


    p138_in <= x(16) & x(20) & x(31) & x(54) & x(138) & x(190) & x(202) & x(208) & x(236) & x(241);
    y(138) <= not(p138_out);
    p138 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1011010000",
            TABLE => "0000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010011110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 5,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p138_in,
            y(0) => p138_out,
            y(1 to 14 - 1) => dummy138
        );


    p139_in <= x(9) & x(30) & x(35) & x(78) & x(113) & x(185) & x(190) & x(208) & x(209);
    y(139) <= not(p139_out);
    p139 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011010011",
            TABLE => "001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p139_in,
            y(0) => p139_out,
            y(1 to 14 - 1) => dummy139
        );


    p140_in <= x(7) & x(8) & x(36) & x(66) & x(69) & x(89) & x(94) & x(125) & x(129) & x(146) & x(149) & x(153) & x(173) & x(179) & x(185) & x(186) & x(207) & x(219) & x(245) & x(247);
    y(140) <= not(p140_out);
    p140 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10011011100111011011",
            TABLE => "001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p140_in,
            y(0) => p140_out,
            y(1 to 14 - 1) => dummy140
        );


    p141_in <= x(9) & x(27) & x(30) & x(36) & x(49) & x(75) & x(78) & x(84) & x(87) & x(89) & x(91) & x(95) & x(101) & x(107) & x(131) & x(137) & x(150) & x(170) & x(174) & x(184) & x(213) & x(222) & x(228) & x(237) & x(244) & x(245);
    y(141) <= not(p141_out);
    p141 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00100101111111000000110111",
            TABLE => "110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p141_in,
            y(0) => p141_out,
            y(1 to 14 - 1) => dummy141
        );


    p142_in <= x(5) & x(6) & x(31) & x(61) & x(82) & x(87) & x(102) & x(103) & x(131) & x(144) & x(154) & x(197) & x(205) & x(206) & x(207) & x(211) & x(241);
    y(142) <= not(p142_out);
    p142 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001001101100101",
            TABLE => "11111011101100101011001000100000101100100010000000100000000000001101101110110010101100100010010010110010001001000010010001001101011010011001011010010110011010011001011001101001011010011001011000010000011100010111000111110111000000000001000000010000011100010001100001110001011100011110011110001110000110000001100001110001100101100110100101101001100101100110100110010110100101100110100111011111010011010100110100000100110110110100110101001101001001001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p142_in,
            y(0) => p142_out,
            y(1 to 14 - 1) => dummy142
        );


    p143_in <= x(34) & x(37) & x(48) & x(57) & x(66) & x(83) & x(102) & x(105) & x(113) & x(121) & x(125) & x(152) & x(185) & x(207) & x(216) & x(224) & x(232) & x(247);
    y(143) <= not(p143_out);
    p143 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100101111101101000",
            TABLE => "010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p143_in,
            y(0) => p143_out,
            y(1 to 14 - 1) => dummy143
        );


    p144_in <= x(5) & x(6) & x(26) & x(29) & x(38) & x(40) & x(47) & x(58) & x(62) & x(70) & x(74) & x(83) & x(112) & x(123) & x(133) & x(138) & x(158) & x(192) & x(221) & x(238) & x(240);
    y(144) <= not(p144_out);
    p144 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111010110110010001010",
            TABLE => "000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001101100101001011011111111",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p144_in,
            y(0) => p144_out,
            y(1 to 14 - 1) => dummy144
        );


    p145_in <= x(4) & x(9) & x(10) & x(31) & x(113) & x(121) & x(126) & x(144) & x(191) & x(208) & x(222) & x(230) & x(243);
    y(145) <= not(p145_out);
    p145 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000111101100",
            TABLE => "1111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010000001000000000001010110000001000101011000000101011111100101011010000101101010000101011010000100010101101000010101111010010101110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 5,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p145_in,
            y(0) => p145_out,
            y(1 to 14 - 1) => dummy145
        );


    p146_in <= x(4) & x(17) & x(28) & x(56) & x(62) & x(84) & x(85) & x(90) & x(115) & x(117) & x(125) & x(132) & x(144) & x(167) & x(174) & x(199) & x(211) & x(213) & x(237) & x(239) & x(246);
    y(146) <= not(p146_out);
    p146 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010110011110001110011",
            TABLE => "001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 4,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p146_in,
            y(0) => p146_out,
            y(1 to 14 - 1) => dummy146
        );


    p147_in <= x(2) & x(6) & x(30) & x(208) & x(220);
    y(147) <= not(p147_out);
    p147 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01000",
            TABLE => "11101000111111101000000011101000111010000111111010000001111010000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 6,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p147_in,
            y(0) => p147_out,
            y(1 to 14 - 1) => dummy147
        );


    p148_in <= x(1) & x(6) & x(8) & x(20) & x(33) & x(38) & x(49) & x(53) & x(57) & x(65) & x(80) & x(83) & x(102) & x(103) & x(118) & x(181) & x(199) & x(211) & x(233);
    y(148) <= not(p148_out);
    p148 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100011100000110001",
            TABLE => "1101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010011000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p148_in,
            y(0) => p148_out,
            y(1 to 14 - 1) => dummy148
        );


    p149_in <= x(14) & x(31) & x(37) & x(44) & x(52) & x(56) & x(60) & x(91) & x(99) & x(112) & x(151) & x(158) & x(192) & x(205) & x(213) & x(223) & x(226) & x(243) & x(248) & x(251);
    y(149) <= not(p149_out);
    p149 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01101110101010010101",
            TABLE => "000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p149_in,
            y(0) => p149_out,
            y(1 to 14 - 1) => dummy149
        );


    p150_in <= x(8) & x(9) & x(14) & x(23) & x(27) & x(30) & x(32) & x(36) & x(61) & x(78) & x(84) & x(95) & x(104) & x(107) & x(115) & x(119) & x(120) & x(125) & x(132) & x(140) & x(148) & x(181) & x(183) & x(222) & x(237) & x(239) & x(245);
    y(150) <= not(p150_out);
    p150 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001101000011110011111011101",
            TABLE => "010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110010011010110100111111111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p150_in,
            y(0) => p150_out,
            y(1 to 14 - 1) => dummy150
        );


    p151_in <= x(40) & x(46) & x(67) & x(68) & x(70) & x(86) & x(97) & x(106) & x(128) & x(131) & x(137) & x(158) & x(164) & x(186) & x(191) & x(192) & x(200) & x(215) & x(227) & x(233) & x(236) & x(240) & x(253);
    y(151) <= not(p151_out);
    p151 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10110000000010101000011",
            TABLE => "00001000100011100000000000001000100011101110111100001000100011100001100010001110011100010001100010001110111001110001100010001110011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000111010001000000010000000000000000111111011101000111010001000000111101000100000011000000100010111100101100110100101101001100101100110100110010110100101100110100100100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011011110111011100010111000100010000111001110111000101110001000110001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p151_in,
            y(0) => p151_out,
            y(1 to 14 - 1) => dummy151
        );


    p152_in <= x(8) & x(23) & x(36) & x(41) & x(85) & x(89) & x(106) & x(125) & x(138) & x(158) & x(164) & x(170) & x(180) & x(184) & x(191) & x(196) & x(213) & x(225) & x(253);
    y(152) <= not(p152_out);
    p152 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0101001111011100000",
            TABLE => "1000111000001000111011111000111000001000000000001000111000001000100011100001100011100111100011100001100001110001100011100001100010010110011010010110100110010110011010011001011010010110011010010000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101101000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p152_in,
            y(0) => p152_out,
            y(1 to 14 - 1) => dummy152
        );


    p153_in <= x(11) & x(41) & x(58) & x(65) & x(75) & x(85) & x(101) & x(105) & x(111) & x(115) & x(142) & x(152) & x(164) & x(176) & x(189) & x(194) & x(201) & x(203) & x(206) & x(232) & x(237) & x(246) & x(247) & x(252);
    y(153) <= not(p153_out);
    p153 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100001001100100100010111",
            TABLE => "110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p153_in,
            y(0) => p153_out,
            y(1 to 14 - 1) => dummy153
        );


    p154_in <= x(17) & x(18) & x(35) & x(46) & x(51) & x(60) & x(64) & x(65) & x(119) & x(127) & x(137) & x(162) & x(164) & x(165) & x(168) & x(186) & x(200) & x(203) & x(205) & x(208) & x(223) & x(235) & x(247);
    y(154) <= not(p154_out);
    p154 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10111001100111111001101",
            TABLE => "00000010001010110000000000000010001010111011111100000010001010110100001000101011110101000100001000101011101111010100001000101011100101100110100101101001100101100110100110010110100101100110100101000000110101001101010011111101000000000100000001000000110101000100001011010100110101001011110100101011010000100100001011010100011010011001011010010110011010011001011001101001011010011001011000000000000000100000001000101011000000100010101100101011101111111101010001000010010000100010101101000010001010110010101110111101011010011001011010010110011010011001011001101001011010011001011001001101110111110000010001001101010011011101101100100100010011010110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p154_in,
            y(0) => p154_out,
            y(1 to 14 - 1) => dummy154
        );


    p155_in <= x(17) & x(27) & x(40) & x(51) & x(56) & x(80) & x(84) & x(86) & x(99) & x(104) & x(128) & x(133) & x(134) & x(135) & x(137) & x(138) & x(139) & x(145) & x(172) & x(177) & x(178) & x(186) & x(215) & x(222) & x(227) & x(233) & x(244) & x(251) & x(253) & x(254);
    y(155) <= not(p155_out);
    p155 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010000010010111011001110110001",
            TABLE => "111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p155_in,
            y(0) => p155_out,
            y(1 to 15 - 1) => dummy155
        );


    p156_in <= x(5) & x(38) & x(74) & x(77) & x(134) & x(138) & x(152) & x(188) & x(196) & x(248);
    y(156) <= not(p156_out);
    p156 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111011101",
            TABLE => "0000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100000010001001101001001000100110110010110011010010000000000000000",
            SHIFT => 5,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p156_in,
            y(0) => p156_out,
            y(1 to 14 - 1) => dummy156
        );


    p157_in <= x(28) & x(29) & x(33) & x(48) & x(52) & x(65) & x(72) & x(88) & x(92) & x(94) & x(97) & x(113) & x(117) & x(135) & x(137) & x(148) & x(155) & x(156) & x(158) & x(170) & x(172) & x(177) & x(200) & x(222) & x(223) & x(251) & x(252) & x(253);
    y(157) <= not(p157_out);
    p157 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101000011100110001100000010",
            TABLE => "0000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101100010101110111111000000100010101100000010001010110000000000000010001010111011110101000010001010110100001000101011110101000100001001101001100101101001011001101001100101100110100101101001100101101000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010011000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011011001000100000101100100010010010010110011010010000000000000000",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p157_in,
            y(0) => p157_out,
            y(1 to 14 - 1) => dummy157
        );


    p158_in <= x(11) & x(27) & x(40) & x(55) & x(65) & x(66) & x(82) & x(90) & x(91) & x(93) & x(96) & x(107) & x(141) & x(150) & x(152) & x(174) & x(186) & x(188) & x(204) & x(240);
    y(158) <= not(p158_out);
    p158 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01011101010011011010",
            TABLE => "000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p158_in,
            y(0) => p158_out,
            y(1 to 14 - 1) => dummy158
        );


    p159_in <= x(4) & x(17) & x(19) & x(21) & x(36) & x(42) & x(60) & x(66) & x(68) & x(88) & x(94) & x(96) & x(115) & x(117) & x(140) & x(167) & x(175) & x(176) & x(180) & x(186) & x(187) & x(197) & x(199) & x(219) & x(223) & x(226) & x(232) & x(237) & x(238) & x(251) & x(254);
    y(159) <= not(p159_out);
    p159 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110001011011100111010111000110",
            TABLE => "1000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010010001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010010001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010010111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p159_in,
            y(0) => p159_out,
            y(1 to 15 - 1) => dummy159
        );


    p160_in <= x(2) & x(5) & x(6) & x(16) & x(19) & x(25) & x(37) & x(57) & x(106) & x(140) & x(141) & x(150) & x(153) & x(181) & x(185) & x(190) & x(207) & x(240) & x(245) & x(248) & x(252);
    y(160) <= not(p160_out);
    p160 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100011100100100011101",
            TABLE => "011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110010011010110100111111111",
            SHIFT => 4,
            B => 8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p160_in,
            y(0) => p160_out,
            y(1 to 14 - 1) => dummy160
        );


    p161_in <= x(7) & x(23) & x(25) & x(48) & x(52) & x(62) & x(76) & x(84) & x(94) & x(96) & x(98) & x(125) & x(135) & x(173) & x(179) & x(220) & x(228) & x(229) & x(233) & x(245);
    y(161) <= not(p161_out);
    p161 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11011110101111101111",
            TABLE => "000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p161_in,
            y(0) => p161_out,
            y(1 to 14 - 1) => dummy161
        );


    p162_in <= x(31) & x(51) & x(64) & x(87) & x(99) & x(110) & x(123) & x(134) & x(151) & x(172) & x(178) & x(202) & x(212) & x(213) & x(230);
    y(162) <= not(p162_out);
    p162 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000100010011110",
            TABLE => "111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110001010110110100111111111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p162_in,
            y(0) => p162_out,
            y(1 to 13 - 1) => dummy162
        );


    p163_in <= x(11) & x(29) & x(36) & x(75) & x(78) & x(93) & x(95) & x(200) & x(201) & x(206) & x(246);
    y(163) <= not(p163_out);
    p163 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101101001",
            TABLE => "01110001111101110001000001110001000100000111000100000000000100000111000111100111000110000111000100011000011100011000111000011000011010011001011010010110011010011001011001101001011010011001011011010100111111010100000011010100110101001011110101000010110101001001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -10,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p163_in,
            y(0) => p163_out,
            y(1 to 13 - 1) => dummy163
        );


    p164_in <= x(8) & x(22) & x(37) & x(42) & x(63) & x(66) & x(73) & x(76) & x(85) & x(129) & x(140) & x(141) & x(146) & x(150) & x(155) & x(159) & x(179) & x(180) & x(188) & x(192) & x(202) & x(225) & x(233) & x(245);
    y(164) <= not(p164_out);
    p164 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011111010110000010010011",
            TABLE => "000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p164_in,
            y(0) => p164_out,
            y(1 to 14 - 1) => dummy164
        );


    p165_in <= x(11) & x(14) & x(15) & x(27) & x(36) & x(40) & x(51) & x(56) & x(59) & x(62) & x(86) & x(99) & x(131) & x(138) & x(145) & x(171) & x(178) & x(186) & x(190) & x(203) & x(215) & x(221) & x(233) & x(240) & x(244);
    y(165) <= not(p165_out);
    p165 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001100000101011110110100",
            TABLE => "1011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p165_in,
            y(0) => p165_out,
            y(1 to 14 - 1) => dummy165
        );


    p166_in <= x(18) & x(35) & x(46) & x(50) & x(51) & x(65) & x(76) & x(90) & x(117) & x(119) & x(134) & x(138) & x(165) & x(168) & x(189) & x(194) & x(235) & x(239) & x(241);
    y(166) <= not(p166_out);
    p166 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0110111111011101011",
            TABLE => "0001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p166_in,
            y(0) => p166_out,
            y(1 to 14 - 1) => dummy166
        );


    p167_in <= x(4) & x(31) & x(35) & x(58) & x(73) & x(76) & x(82) & x(123) & x(130) & x(140) & x(142) & x(146) & x(168) & x(170) & x(175) & x(191) & x(196) & x(202) & x(211) & x(236) & x(249);
    y(167) <= not(p167_out);
    p167 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "000010000001011001110",
            TABLE => "111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110001010110110100111111111",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p167_in,
            y(0) => p167_out,
            y(1 to 14 - 1) => dummy167
        );


    p168_in <= x(13) & x(52) & x(60) & x(73) & x(89) & x(90) & x(93) & x(115) & x(117) & x(125) & x(149) & x(152) & x(167) & x(175) & x(182) & x(197) & x(224) & x(234) & x(251) & x(253);
    y(168) <= not(p168_out);
    p168 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10001000001110111000",
            TABLE => "101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p168_in,
            y(0) => p168_out,
            y(1 to 14 - 1) => dummy168
        );


    p169_in <= x(11) & x(22) & x(28) & x(37) & x(46) & x(56) & x(65) & x(84) & x(86) & x(105) & x(106) & x(110) & x(140) & x(146) & x(191) & x(202) & x(211) & x(228) & x(232) & x(236) & x(239) & x(240);
    y(169) <= not(p169_out);
    p169 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100101011100101110110",
            TABLE => "1011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010010000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010010010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p169_in,
            y(0) => p169_out,
            y(1 to 14 - 1) => dummy169
        );


    p170_in <= x(2) & x(40) & x(46) & x(68) & x(78) & x(86) & x(96) & x(97) & x(128) & x(135) & x(137) & x(150) & x(170) & x(177) & x(186) & x(191) & x(222) & x(227) & x(240) & x(244) & x(253) & x(254);
    y(170) <= not(p170_out);
    p170 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101001000000101101110",
            TABLE => "0000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101101110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101100010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101100000001000101011010000100010101110010110011010010000000000000000",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p170_in,
            y(0) => p170_out,
            y(1 to 14 - 1) => dummy170
        );


    p171_in <= x(2) & x(9) & x(15) & x(16) & x(24) & x(55) & x(64) & x(68) & x(74) & x(80) & x(87) & x(94) & x(119) & x(142) & x(144) & x(154) & x(158) & x(183) & x(238) & x(253);
    y(171) <= not(p171_out);
    p171 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10100111110000010111",
            TABLE => "010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001000110010000",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p171_in,
            y(0) => p171_out,
            y(1 to 14 - 1) => dummy171
        );


    p172_in <= x(3) & x(11) & x(17) & x(28) & x(32) & x(51) & x(65) & x(77) & x(120) & x(127) & x(129) & x(137) & x(157) & x(158) & x(164) & x(165) & x(168) & x(173) & x(193) & x(205) & x(219) & x(223) & x(230) & x(239) & x(241);
    y(172) <= not(p172_out);
    p172 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101000011110100010100000",
            TABLE => "0000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101100001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010011101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010011110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p172_in,
            y(0) => p172_out,
            y(1 to 14 - 1) => dummy172
        );


    p173_in <= x(1) & x(17) & x(28) & x(32) & x(33) & x(37) & x(51) & x(62) & x(65) & x(87) & x(88) & x(90) & x(167) & x(185) & x(187) & x(193) & x(199) & x(204) & x(232) & x(236) & x(249);
    y(173) <= not(p173_out);
    p173 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110110101011011111010",
            TABLE => "000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => 4,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p173_in,
            y(0) => p173_out,
            y(1 to 14 - 1) => dummy173
        );


    p174_in <= x(1) & x(58) & x(65) & x(83) & x(116) & x(118) & x(120) & x(134) & x(138) & x(147) & x(170) & x(181) & x(197) & x(207) & x(224) & x(235);
    y(174) <= not(p174_out);
    p174 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1011100011110000",
            TABLE => "0000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010011110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p174_in,
            y(0) => p174_out,
            y(1 to 14 - 1) => dummy174
        );


    p175_in <= x(15) & x(36) & x(44) & x(48) & x(52) & x(59) & x(87) & x(89) & x(130) & x(155) & x(174) & x(175) & x(179) & x(180) & x(200) & x(216) & x(224) & x(226) & x(238) & x(252) & x(253);
    y(175) <= not(p175_out);
    p175 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011100111000000111010",
            TABLE => "000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p175_in,
            y(0) => p175_out,
            y(1 to 14 - 1) => dummy175
        );


    p176_in <= x(7) & x(14) & x(18) & x(19) & x(32) & x(38) & x(52) & x(55) & x(62) & x(67) & x(74) & x(84) & x(93) & x(125) & x(135) & x(153) & x(159) & x(164) & x(172) & x(173) & x(233) & x(245);
    y(176) <= not(p176_out);
    p176 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110011111101111011111",
            TABLE => "0000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010010000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100000000100010111100000010001011101101001100101100000000000000000",
            SHIFT => 4,
            B => -6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p176_in,
            y(0) => p176_out,
            y(1 to 14 - 1) => dummy176
        );


    p177_in <= x(14) & x(24) & x(32) & x(37) & x(48) & x(71) & x(85) & x(91) & x(94) & x(96) & x(97) & x(113) & x(121) & x(136) & x(146) & x(184) & x(186) & x(187) & x(213) & x(222) & x(233) & x(243);
    y(177) <= not(p177_out);
    p177 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1000001101011110011100",
            TABLE => "1110100010000000100000000000000011111110111010001110100010000000111010001000000110000001000101110111111011101000111010001000000101101001100101101001011001101001100101100110100101101001100101100000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010010000100010001110000110001000111001101001100101100000000000000000",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p177_in,
            y(0) => p177_out,
            y(1 to 14 - 1) => dummy177
        );


    p178_in <= x(18) & x(52) & x(59) & x(84) & x(94) & x(102) & x(148) & x(157) & x(162) & x(172) & x(173) & x(177) & x(216) & x(221) & x(229) & x(237) & x(250) & x(253) & x(254);
    y(178) <= not(p178_out);
    p178 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001100110001001101",
            TABLE => "1011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p178_in,
            y(0) => p178_out,
            y(1 to 14 - 1) => dummy178
        );


    p179_in <= x(5) & x(17) & x(43) & x(51) & x(56) & x(92) & x(93) & x(99) & x(111) & x(127) & x(134) & x(135) & x(138) & x(147) & x(182) & x(194) & x(207) & x(213) & x(218) & x(225) & x(232) & x(241) & x(244) & x(251);
    y(179) <= not(p179_out);
    p179 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010111011000111100111111",
            TABLE => "000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p179_in,
            y(0) => p179_out,
            y(1 to 14 - 1) => dummy179
        );


    p180_in <= x(14) & x(17) & x(26) & x(51) & x(63) & x(74) & x(91) & x(100) & x(107) & x(116) & x(126) & x(137) & x(144) & x(149) & x(162) & x(203) & x(229) & x(237);
    y(180) <= not(p180_out);
    p180 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110100101110101001",
            TABLE => "000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 5,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p180_in,
            y(0) => p180_out,
            y(1 to 15 - 1) => dummy180
        );


    p181_in <= x(8) & x(14) & x(16) & x(27) & x(30) & x(32) & x(70) & x(80) & x(87) & x(91) & x(95) & x(103) & x(107) & x(117) & x(118) & x(123) & x(125) & x(126) & x(132) & x(136) & x(143) & x(186) & x(192) & x(201) & x(218) & x(222) & x(230) & x(245);
    y(181) <= not(p181_out);
    p181 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100100111111010111100011101",
            TABLE => "1011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010010000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100001000001110001000000000001000001110001111101110001000001110001000110000111000110001110000110000111000111100111000110000111000110010110011010010110100110010110011010011001011010010110011010010100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101100000010001001101001001000100110110010110011010010000000000000000",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p181_in,
            y(0) => p181_out,
            y(1 to 14 - 1) => dummy181
        );


    p182_in <= x(5) & x(6) & x(30) & x(57) & x(76) & x(81) & x(96) & x(121) & x(123) & x(138) & x(198) & x(199) & x(202) & x(205) & x(212) & x(238);
    y(182) <= not(p182_out);
    p182 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101110010000101",
            TABLE => "0000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101101110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100100110100000100010011010010010001101001100101100000000000000000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p182_in,
            y(0) => p182_out,
            y(1 to 14 - 1) => dummy182
        );


    p183_in <= x(14) & x(32) & x(50) & x(62) & x(82) & x(87) & x(91) & x(112) & x(116) & x(151) & x(171) & x(192) & x(213) & x(224) & x(241);
    y(183) <= not(p183_out);
    p183 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011000000111011",
            TABLE => "100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110011100010110100111111111",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p183_in,
            y(0) => p183_out,
            y(1 to 13 - 1) => dummy183
        );


    p184_in <= x(2) & x(9) & x(24) & x(27) & x(67) & x(68) & x(94) & x(97) & x(119) & x(120) & x(121) & x(124) & x(154) & x(158) & x(170) & x(177) & x(185) & x(186) & x(220) & x(222) & x(227) & x(231) & x(238) & x(247) & x(253) & x(254);
    y(184) <= not(p184_out);
    p184 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10001100011110010011001010",
            TABLE => "011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p184_in,
            y(0) => p184_out,
            y(1 to 14 - 1) => dummy184
        );


    p185_in <= x(25) & x(38) & x(48) & x(66) & x(85) & x(98) & x(122) & x(137) & x(153) & x(162) & x(163) & x(173) & x(185) & x(208) & x(209) & x(214) & x(220) & x(230) & x(231) & x(239);
    y(185) <= not(p185_out);
    p185 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110010010001100101",
            TABLE => "000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110010001100000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p185_in,
            y(0) => p185_out,
            y(1 to 14 - 1) => dummy185
        );


    p186_in <= x(10) & x(14) & x(32) & x(37) & x(53) & x(82) & x(84) & x(102) & x(110) & x(116) & x(141) & x(151) & x(175) & x(192) & x(196) & x(213) & x(219) & x(224) & x(241);
    y(186) <= not(p186_out);
    p186 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1011101010010100111",
            TABLE => "0000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p186_in,
            y(0) => p186_out,
            y(1 to 14 - 1) => dummy186
        );


    p187_in <= x(4) & x(5) & x(14) & x(20) & x(26) & x(36) & x(50) & x(52) & x(57) & x(60) & x(67) & x(72) & x(98) & x(102) & x(110) & x(112) & x(125) & x(151) & x(170) & x(190) & x(191) & x(192) & x(213) & x(219) & x(223) & x(226) & x(251);
    y(187) <= not(p187_out);
    p187 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111101001001110100110010010",
            TABLE => "000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p187_in,
            y(0) => p187_out,
            y(1 to 14 - 1) => dummy187
        );


    p188_in <= x(11) & x(20) & x(22) & x(29) & x(79) & x(82) & x(93) & x(137) & x(165) & x(176) & x(179) & x(180) & x(200) & x(213) & x(253);
    y(188) <= not(p188_out);
    p188 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100110010101000",
            TABLE => "001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p188_in,
            y(0) => p188_out,
            y(1 to 13 - 1) => dummy188
        );


    p189_in <= x(5) & x(11) & x(22) & x(25) & x(29) & x(47) & x(56) & x(70) & x(99) & x(113) & x(117) & x(126) & x(141) & x(246);
    y(189) <= not(p189_out);
    p189 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10100101011011",
            TABLE => "010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 5,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p189_in,
            y(0) => p189_out,
            y(1 to 14 - 1) => dummy189
        );


    p190_in <= x(8) & x(17) & x(31) & x(35) & x(36) & x(43) & x(75) & x(85) & x(95) & x(103) & x(125) & x(138) & x(152) & x(158) & x(196) & x(200) & x(219) & x(253);
    y(190) <= not(p190_out);
    p190 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010000101111110000",
            TABLE => "111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p190_in,
            y(0) => p190_out,
            y(1 to 14 - 1) => dummy190
        );


    p191_in <= x(125) & x(135) & x(162) & x(208) & x(210) & x(247) & x(250);
    y(191) <= not(p191_out);
    p191 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111011",
            TABLE => "0000000000000100000001000100110100000100010011010100110111011111101100100010010000100100010011010010010001001101010011011101101101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p191_in,
            y(0) => p191_out,
            y(1 to 13 - 1) => dummy191
        );


    p192_in <= x(15) & x(48) & x(53) & x(58) & x(72) & x(73) & x(84) & x(114) & x(138) & x(155) & x(167) & x(203) & x(219) & x(252);
    y(192) <= not(p192_out);
    p192 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110010001111",
            TABLE => "000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p192_in,
            y(0) => p192_out,
            y(1 to 13 - 1) => dummy192
        );


    p193_in <= x(3) & x(8) & x(29) & x(62) & x(89) & x(94) & x(95) & x(123) & x(125) & x(126) & x(138) & x(168) & x(170) & x(181) & x(184) & x(201) & x(208) & x(217) & x(218) & x(230) & x(246) & x(249) & x(253);
    y(193) <= not(p193_out);
    p193 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10110110111010111010000",
            TABLE => "00000100010011010000000000000100010011011101111100000100010011010010010001001101101100100010010001001101110110110010010001001101100101100110100101101001100101100110100110010110100101100110100100000010001010110000000000000010001010111011111100000010001010110100001000101011110101000100001000101011101111010100001000101011100101100110100101101001100101100110100110010110100101100110100100000010001010110000000000000010001010111011111100000010001010110100001000101011110101000100001000101011101111010100001000101011100101100110100101101001100101100110100110010110100101100110100111101000100000001111111011101000111010001000000101111110111010000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p193_in,
            y(0) => p193_out,
            y(1 to 14 - 1) => dummy193
        );


    p194_in <= x(9) & x(20) & x(21) & x(29) & x(60) & x(69) & x(74) & x(97) & x(100) & x(111) & x(117) & x(132) & x(134) & x(147) & x(150) & x(162) & x(180) & x(194) & x(206) & x(208) & x(237) & x(238) & x(248) & x(250) & x(253);
    y(194) <= not(p194_out);
    p194 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001101111100110111001000",
            TABLE => "0010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010011000111000001000000010000000000011101111100011101000111000001000100011100001100000011000011100011110011110001110100011100001100010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p194_in,
            y(0) => p194_out,
            y(1 to 14 - 1) => dummy194
        );


    p195_in <= x(1) & x(6) & x(24) & x(66) & x(91) & x(96) & x(105) & x(107) & x(158) & x(163) & x(179) & x(200) & x(204) & x(205) & x(206) & x(213) & x(253);
    y(195) <= not(p195_out);
    p195 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001111110000110",
            TABLE => "11110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100100000000000010000000100010001110000010001000111010001110111011110111000100011000000110001000111000011000100011101000111011100111100101100110100101101001100101100110100110010110100101100110100110111111001010110010101100000010101111010010101100101011010000101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p195_in,
            y(0) => p195_out,
            y(1 to 14 - 1) => dummy195
        );


    p196_in <= x(36) & x(50) & x(52) & x(56) & x(70) & x(82) & x(88) & x(112) & x(153) & x(154) & x(164) & x(165) & x(168) & x(175) & x(176) & x(203) & x(207) & x(210) & x(232) & x(240) & x(244) & x(245) & x(247);
    y(196) <= not(p196_out);
    p196 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00110101101110000011111",
            TABLE => "01001101110111110000010001001101000001000100110100000000000001000100110111011011001001000100110100100100010011011011001000100100011010011001011010010110011010011001011001101001011010011001011000010000011100010111000111110111000000000001000000010000011100010001100001110001011100011110011110001110000110000001100001110001100101100110100101101001100101100110100110010110100101100110100111101000100000001000000000000000111111101110100011101000100000001110100010000001100000010001011101111110111010001110100010000001011010011001011010010110011010011001011001101001011010011001011000000001000101110001011101111111100000010001011100010111011111100110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p196_in,
            y(0) => p196_out,
            y(1 to 14 - 1) => dummy196
        );


    p197_in <= x(63) & x(85) & x(225) & x(228) & x(247);
    y(197) <= not(p197_out);
    p197 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110",
            TABLE => "00101011101111110000001000101011001010111011110101000010001010110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 6,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p197_in,
            y(0) => p197_out,
            y(1 to 14 - 1) => dummy197
        );


    p198_in <= x(18) & x(19) & x(28) & x(41) & x(65) & x(87) & x(88) & x(99) & x(126) & x(157) & x(158) & x(174) & x(195) & x(208) & x(212) & x(245);
    y(198) <= not(p198_out);
    p198 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010010000100011",
            TABLE => "0100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101101111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100111000100010000011100010001100001101001100101100000000000000000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p198_in,
            y(0) => p198_out,
            y(1 to 14 - 1) => dummy198
        );


    p199_in <= x(7) & x(11) & x(34) & x(38) & x(52) & x(55) & x(65) & x(74) & x(75) & x(83) & x(84) & x(89) & x(90) & x(91) & x(107) & x(116) & x(117) & x(125) & x(132) & x(134) & x(144) & x(145) & x(147) & x(172) & x(192) & x(205) & x(213) & x(216) & x(229) & x(237) & x(239) & x(246) & x(249);
    y(199) <= not(p199_out);
    p199 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100111110000100011000011100010110",
            TABLE => "000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001001010110110100111111111",
            SHIFT => 3,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p199_in,
            y(0) => p199_out,
            y(1 to 14 - 1) => dummy199
        );


    p200_in <= x(2) & x(18) & x(26) & x(41) & x(67) & x(94) & x(101) & x(103) & x(132) & x(160) & x(162) & x(170) & x(172) & x(177) & x(186) & x(191) & x(195) & x(208) & x(241) & x(250) & x(254);
    y(200) <= not(p200_out);
    p200 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "111010100100110100000",
            TABLE => "000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p200_in,
            y(0) => p200_out,
            y(1 to 14 - 1) => dummy200
        );


    p201_in <= x(10) & x(14) & x(37) & x(39) & x(41) & x(63) & x(69) & x(76) & x(83) & x(102) & x(103) & x(108) & x(109) & x(113) & x(121) & x(131) & x(132) & x(161) & x(162) & x(184) & x(185) & x(192) & x(196) & x(199) & x(206) & x(212) & x(255);
    y(201) <= not(p201_out);
    p201 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101010100010000110110100000",
            TABLE => "001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p201_in,
            y(0) => p201_out,
            y(1 to 14 - 1) => dummy201
        );


    p202_in <= x(18) & x(48) & x(63) & x(66) & x(89) & x(113) & x(122) & x(123) & x(134) & x(137) & x(144) & x(149) & x(158) & x(162) & x(164) & x(173) & x(194) & x(207) & x(214) & x(216) & x(220) & x(230) & x(231) & x(252);
    y(202) <= not(p202_out);
    p202 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "101000001101100101101010",
            TABLE => "100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p202_in,
            y(0) => p202_out,
            y(1 to 14 - 1) => dummy202
        );


    p203_in <= x(18) & x(26) & x(38) & x(47) & x(49) & x(56) & x(58) & x(59) & x(62) & x(66) & x(67) & x(74) & x(80) & x(99) & x(123) & x(126) & x(142) & x(170) & x(216) & x(221) & x(241) & x(244);
    y(203) <= not(p203_out);
    p203 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111101001110010100000",
            TABLE => "0000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010011011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010011110100010000000111010001000000101101001100101100000000000000000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p203_in,
            y(0) => p203_out,
            y(1 to 14 - 1) => dummy203
        );


    p204_in <= x(85) & x(96) & x(152) & x(157) & x(198) & x(203) & x(206) & x(226);
    y(204) <= not(p204_out);
    p204 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01101110",
            TABLE => "000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001001001100000",
            SHIFT => 5,
            B => -9,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p204_in,
            y(0) => p204_out,
            y(1 to 14 - 1) => dummy204
        );


    p205_in <= x(10) & x(15) & x(83) & x(102) & x(105) & x(109) & x(113) & x(119) & x(120) & x(127) & x(129) & x(143) & x(152) & x(179) & x(182) & x(193) & x(203) & x(225);
    y(205) <= not(p205_out);
    p205 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001111110001101101",
            TABLE => "000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p205_in,
            y(0) => p205_out,
            y(1 to 14 - 1) => dummy205
        );


    p206_in <= x(4) & x(61) & x(87) & x(99) & x(110) & x(116) & x(117) & x(123) & x(144) & x(147) & x(179) & x(200) & x(206) & x(212) & x(230) & x(247) & x(253);
    y(206) <= not(p206_out);
    p206 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01100100100011000",
            TABLE => "01000000110101001101010011111101000000000100000001000000110101000100001011010100110101001011110100101011010000100100001011010100011010011001011010010110011010011001011001101001011010011001011011101000111111101000000011101000100000001110100000000000100000001110100001111110100000011110100010000001111010000001011110000001011010011001011010010110011010011001011001101001011010011001011010000000111010001110100011111110100000011110100011101000011111101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p206_in,
            y(0) => p206_out,
            y(1 to 14 - 1) => dummy206
        );


    p207_in <= x(6) & x(14) & x(16) & x(29) & x(32) & x(36) & x(65) & x(91) & x(118) & x(123) & x(152) & x(158) & x(171) & x(173) & x(183) & x(185) & x(195) & x(200) & x(230) & x(239) & x(243);
    y(207) <= not(p207_out);
    p207 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010100011011111000000",
            TABLE => "100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110111010000110100111111111",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p207_in,
            y(0) => p207_out,
            y(1 to 14 - 1) => dummy207
        );


    p208_in <= x(5) & x(6) & x(16) & x(32) & x(48) & x(49) & x(87) & x(91) & x(99) & x(107) & x(112) & x(116) & x(151) & x(152) & x(161) & x(190) & x(195) & x(236) & x(241);
    y(208) <= not(p208_out);
    p208 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001100010001110111",
            TABLE => "1011111100101011001010110000001000101011000000100000001000000000101111010010101100101011010000100010101101000010010000101101010010010110011010010110100110010110011010011001011010010110011010011110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p208_in,
            y(0) => p208_out,
            y(1 to 14 - 1) => dummy208
        );


    p209_in <= x(0) & x(7) & x(32) & x(35) & x(36) & x(60) & x(79) & x(122) & x(129) & x(140) & x(146) & x(153) & x(154) & x(173) & x(180) & x(193) & x(196) & x(213) & x(235) & x(237) & x(238) & x(245) & x(247) & x(249);
    y(209) <= not(p209_out);
    p209 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110100011101010011010111",
            TABLE => "000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p209_in,
            y(0) => p209_out,
            y(1 to 14 - 1) => dummy209
        );


    p210_in <= x(8) & x(21) & x(35) & x(40) & x(70) & x(84) & x(86) & x(87) & x(97) & x(101) & x(107) & x(115) & x(117) & x(118) & x(132) & x(175) & x(180) & x(194) & x(196) & x(211) & x(213) & x(234) & x(237) & x(238) & x(240) & x(245);
    y(210) <= not(p210_out);
    p210 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01110101011001100010101011",
            TABLE => "000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110000110010000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p210_in,
            y(0) => p210_out,
            y(1 to 14 - 1) => dummy210
        );


    p211_in <= x(56) & x(93) & x(99) & x(138) & x(158) & x(171) & x(206);
    y(211) <= not(p211_out);
    p211 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1011101",
            TABLE => "0000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 6,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p211_in,
            y(0) => p211_out,
            y(1 to 14 - 1) => dummy211
        );


    p212_in <= x(2) & x(3) & x(5) & x(6) & x(61) & x(80) & x(102) & x(113) & x(119) & x(121) & x(140) & x(141) & x(144) & x(150) & x(151) & x(163) & x(169) & x(172) & x(177) & x(202) & x(206);
    y(212) <= not(p212_out);
    p212 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011110101001110100001",
            TABLE => "000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110110101001001011011111111",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p212_in,
            y(0) => p212_out,
            y(1 to 14 - 1) => dummy212
        );


    p213_in <= x(24) & x(32) & x(35) & x(40) & x(44) & x(47) & x(51) & x(52) & x(58) & x(62) & x(71) & x(82) & x(89) & x(99) & x(107) & x(110) & x(125) & x(129) & x(143) & x(146) & x(152) & x(196) & x(215) & x(221) & x(238) & x(240) & x(244) & x(251);
    y(213) <= not(p213_out);
    p213 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1011001101110101110001010111",
            TABLE => "0000100010001110000000000000100010001110111011110000100010001110000110001000111001110001000110001000111011100111000110001000111001101001100101101001011001101001100101100110100101101001100101100000000100000000000101110000000100010111000000010111111100010111100000011110100000010111100000010001011110000001011111100001011101101001100101101001011001101001100101100110100101101001100101100001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010011101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010010001011100000001000101111000000110010110011010010000000000000000",
            SHIFT => 3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p213_in,
            y(0) => p213_out,
            y(1 to 13 - 1) => dummy213
        );


    p214_in <= x(8) & x(13) & x(14) & x(34) & x(58) & x(83) & x(85) & x(101) & x(142) & x(153) & x(171) & x(175) & x(189) & x(203) & x(229) & x(233) & x(237) & x(238) & x(245);
    y(214) <= not(p214_out);
    p214 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0100100111101111101",
            TABLE => "1011001000100000111110111011001000100000000000001011001000100000101100100010010011011011101100100010010001001101101100100010010010010110011010010110100110010110011010011001011010010110011010010000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010010000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 5,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p214_in,
            y(0) => p214_out,
            y(1 to 15 - 1) => dummy214
        );


    p215_in <= x(4) & x(10) & x(12) & x(25) & x(30) & x(36) & x(38) & x(41) & x(58) & x(64) & x(85) & x(113) & x(118) & x(121) & x(152) & x(157) & x(171) & x(174) & x(188) & x(237) & x(248);
    y(215) <= not(p215_out);
    p215 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001010111101111010111",
            TABLE => "101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p215_in,
            y(0) => p215_out,
            y(1 to 14 - 1) => dummy215
        );


    p216_in <= x(45) & x(48) & x(67) & x(97) & x(116) & x(135) & x(152) & x(194) & x(253);
    y(216) <= not(p216_out);
    p216 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "001000101",
            TABLE => "111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110010011010110100111111111",
            SHIFT => 5,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p216_in,
            y(0) => p216_out,
            y(1 to 14 - 1) => dummy216
        );


    p217_in <= x(12) & x(23) & x(24) & x(34) & x(52) & x(58) & x(59) & x(62) & x(75) & x(89) & x(101) & x(107) & x(113) & x(123) & x(138) & x(144) & x(147) & x(152) & x(153) & x(170) & x(192) & x(195) & x(204) & x(213) & x(238) & x(251);
    y(217) <= not(p217_out);
    p217 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10010100111111010100000110",
            TABLE => "010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110001001100000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p217_in,
            y(0) => p217_out,
            y(1 to 14 - 1) => dummy217
        );


    p218_in <= x(32) & x(45) & x(58) & x(59) & x(87) & x(91) & x(101) & x(113) & x(119) & x(126) & x(142) & x(147) & x(174) & x(195) & x(213) & x(241) & x(255);
    y(218) <= not(p218_out);
    p218 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10010000010111010",
            TABLE => "10001110000010000000100000000000111011111000111010001110000010001000111000011000000110000111000111100111100011101000111000011000100101100110100101101001100101100110100110010110100101100110100111011111010011010100110100000100010011010000010000000100000000001101101101001101010011010010010001001101001001000010010010110010100101100110100101101001100101100110100110010110100101100110100100100000101100101011001011111011001001001011001010110010110110110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p218_in,
            y(0) => p218_out,
            y(1 to 14 - 1) => dummy218
        );


    p219_in <= x(10) & x(13) & x(14) & x(69) & x(89) & x(93) & x(105) & x(113) & x(125) & x(130) & x(135) & x(143) & x(148) & x(158) & x(170) & x(173) & x(174) & x(176) & x(179) & x(182) & x(186) & x(192) & x(207) & x(210) & x(219) & x(239) & x(247) & x(254);
    y(219) <= not(p219_out);
    p219 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1011010010101111101011100011",
            TABLE => "0000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010011011001011111011001000001011001000100000101100100000000000100000101100101101101100100100101100100010010010110010010011010010010010010110011010010110100110010110011010011001011010010110011010010000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010111000100010000011100010001100001101001100101100000000000000000",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p219_in,
            y(0) => p219_out,
            y(1 to 14 - 1) => dummy219
        );


    p220_in <= x(8) & x(22) & x(27) & x(36) & x(52) & x(84) & x(86) & x(103) & x(118) & x(120) & x(125) & x(126) & x(128) & x(132) & x(143) & x(181) & x(186) & x(219) & x(223) & x(227) & x(228) & x(232) & x(240) & x(244) & x(251);
    y(220) <= not(p220_out);
    p220 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000110111110100011001111",
            TABLE => "1111011101110001011100010001000001110001000100000001000000000000111001110111000101110001000110000111000100011000000110001000111010010110011010010110100110010110011010011001011010010110011010010000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101101101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p220_in,
            y(0) => p220_out,
            y(1 to 14 - 1) => dummy220
        );


    p221_in <= x(5) & x(14) & x(37) & x(40) & x(45) & x(50) & x(58) & x(62) & x(68) & x(74) & x(80) & x(83) & x(85) & x(109) & x(112) & x(116) & x(133) & x(139) & x(142) & x(171) & x(187) & x(192) & x(202) & x(203) & x(207) & x(233) & x(240);
    y(221) <= not(p221_out);
    p221 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010110011011111110001010001",
            TABLE => "001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001110101001001011011111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p221_in,
            y(0) => p221_out,
            y(1 to 14 - 1) => dummy221
        );


    p222_in <= x(9) & x(11) & x(14) & x(16) & x(22) & x(23) & x(27) & x(29) & x(40) & x(73) & x(75) & x(97) & x(120) & x(126) & x(142) & x(177) & x(179) & x(186) & x(222) & x(249) & x(253);
    y(222) <= not(p222_out);
    p222 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100110100001001011010",
            TABLE => "001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p222_in,
            y(0) => p222_out,
            y(1 to 14 - 1) => dummy222
        );


    p223_in <= x(2) & x(18) & x(20) & x(26) & x(32) & x(65) & x(67) & x(74) & x(85) & x(87) & x(101) & x(153) & x(162) & x(170) & x(183) & x(208) & x(216) & x(232) & x(241) & x(243) & x(247) & x(253);
    y(223) <= not(p223_out);
    p223 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1101001111110010010001",
            TABLE => "0000100000000000100011100000100010001110000010001110111110001110000110000111000110001110000110001000111000011000111001111000111001101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010011101010011111101010000001101010001000000110101000000000001000000110101001011110101000010110101000100001011010100001010110100001010010110011010010110100110010110011010011001011010010110011010011101010001000000110101000100001010010110011010010000000000000000",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p223_in,
            y(0) => p223_out,
            y(1 to 14 - 1) => dummy223
        );


    p224_in <= x(15) & x(28) & x(48) & x(52) & x(53) & x(58) & x(61) & x(67) & x(72) & x(89) & x(107) & x(117) & x(126) & x(127) & x(130) & x(167) & x(175) & x(200) & x(223) & x(224) & x(237) & x(251) & x(253);
    y(224) <= not(p224_out);
    p224 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01101100011000110001100",
            TABLE => "00010000011100010111000111110111000000000001000000010000011100010001100001110001011100011110011110001110000110000001100001110001100101100110100101101001100101100110100110010110100101100110100110111111001010110010101100000010001010110000001000000010000000001011110100101011001010110100001000101011010000100100001011010100100101100110100101101001100101100110100110010110100101100110100110001110111011110000100010001110000010001000111000000000000010001000111011100111000110001000111000011000100011100111000100011000100101100110100101101001100101100110100110010110100101100110100110001110111011110000100010001110100011101110011100011000100011101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p224_in,
            y(0) => p224_out,
            y(1 to 14 - 1) => dummy224
        );


    p225_in <= x(1) & x(3) & x(8) & x(24) & x(38) & x(58) & x(63) & x(64) & x(83) & x(102) & x(103) & x(109) & x(118) & x(123) & x(131) & x(154) & x(171) & x(185) & x(199) & x(221) & x(233) & x(248) & x(255);
    y(225) <= not(p225_out);
    p225 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00001101001011111000110",
            TABLE => "11110111011100010111000100010000011100010001000000010000000000001110011101110001011100010001100001110001000110000001100010001110100101100110100101101001100101100110100110010110100101100110100110110010001000001111101110110010001000000000000010110010001000001011001000100100110110111011001000100100010011011011001000100100100101100110100101101001100101100110100110010110100101100110100100000000000000100000001000101011000000100010101100101011101111111101010001000010010000100010101101000010001010110010101110111101011010011001011010010110011010011001011001101001011010011001011010111111001010110010101100000010101111010010101100101011010000101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p225_in,
            y(0) => p225_out,
            y(1 to 14 - 1) => dummy225
        );


    p226_in <= x(14) & x(29) & x(34) & x(43) & x(44) & x(57) & x(89) & x(91) & x(107) & x(112) & x(116) & x(122) & x(123) & x(136) & x(145) & x(153) & x(217) & x(226) & x(230) & x(248);
    y(226) <= not(p226_out);
    p226 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01000000000000010000",
            TABLE => "111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p226_in,
            y(0) => p226_out,
            y(1 to 14 - 1) => dummy226
        );


    p227_in <= x(26) & x(30) & x(36) & x(38) & x(47) & x(62) & x(64) & x(83) & x(96) & x(119) & x(123) & x(159) & x(170) & x(183) & x(216) & x(226) & x(255);
    y(227) <= not(p227_out);
    p227 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11011010101001000",
            TABLE => "00000010000000000010101100000010001010110000001010111111001010110100001011010100001010110100001000101011010000101011110100101011100101100110100101101001100101100110100110010110100101100110100100100000101100100000000000100000101100101111101100100000101100100010010010110010010011010010010010110010110110110010010010110010011010011001011010010110011010011001011001101001011010011001011011101000111111101000000011101000111010000111111010000001111010000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p227_in,
            y(0) => p227_out,
            y(1 to 14 - 1) => dummy227
        );


    p228_in <= x(3) & x(5) & x(6) & x(24) & x(28) & x(32) & x(61) & x(65) & x(68) & x(77) & x(80) & x(87) & x(88) & x(119) & x(131) & x(142) & x(144) & x(154) & x(157) & x(158) & x(172) & x(204) & x(230) & x(239) & x(255);
    y(228) <= not(p228_out);
    p228 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1111101000010101100100001",
            TABLE => "0000000000000010000000100010101100000010001010110010101110111111110101000100001001000010001010110100001000101011001010111011110101101001100101101001011001101001100101100110100101101001100101101101010001000000010000000000000011111101110101001101010001000000110101000100001001000010001010111011110111010100110101000100001010010110011010010110100110010110011010011001011010010110011010010010101100000010101111110010101100000010000000000010101100000010001010110100001010111101001010110100001011010100001010110100001001101001100101101001011001101001100101100110100101101001100101101110100010000000111111101110100010000000000000001110100010000000111010001000000101111110111010001000000100010111111010001000000101101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p228_in,
            y(0) => p228_out,
            y(1 to 14 - 1) => dummy228
        );


    p229_in <= x(2) & x(9) & x(70) & x(94) & x(100) & x(220) & x(240);
    y(229) <= not(p229_out);
    p229 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010011",
            TABLE => "0100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 5,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p229_in,
            y(0) => p229_out,
            y(1 to 13 - 1) => dummy229
        );


    p230_in <= x(14) & x(19) & x(45) & x(50) & x(75) & x(88) & x(94) & x(126) & x(135) & x(158) & x(169) & x(176) & x(178) & x(180) & x(195) & x(198) & x(212) & x(232) & x(255);
    y(230) <= not(p230_out);
    p230 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010001011001000111",
            TABLE => "1000000011101000000000001000000011101000111111101000000011101000100000011110100000010111100000011110100001111110100000011110100010010110011010010110100110010110011010011001011010010110011010010000100010001110000000000000100010001110111011110000100010001110000110001000111001110001000110001000111011100111000110001000111001101001100101101001011001101001100101100110100101101001100101100111000100010000000100000000000011110111011100010111000100010000011100010001100000011000100011101110011101110001011100010001100001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p230_in,
            y(0) => p230_out,
            y(1 to 14 - 1) => dummy230
        );


    p231_in <= x(21) & x(29) & x(36) & x(38) & x(43) & x(69) & x(84) & x(85) & x(93) & x(123) & x(145) & x(163) & x(186) & x(228) & x(251);
    y(231) <= not(p231_out);
    p231 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "010000110001001",
            TABLE => "111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110110101001001011011111111",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p231_in,
            y(0) => p231_out,
            y(1 to 13 - 1) => dummy231
        );


    p232_in <= x(35) & x(50) & x(96) & x(112) & x(116) & x(203) & x(226);
    y(232) <= not(p232_out);
    p232 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1001101",
            TABLE => "0010101100000010000000100000000010111111001010110010101100000010001010110100001001000010110101001011110100101011001010110100001001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 5,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p232_in,
            y(0) => p232_out,
            y(1 to 13 - 1) => dummy232
        );


    p233_in <= x(1) & x(20) & x(28) & x(65) & x(85) & x(106) & x(127) & x(134) & x(143) & x(162) & x(173) & x(175) & x(182) & x(189) & x(194) & x(209) & x(231) & x(235) & x(239) & x(247);
    y(233) <= not(p233_out);
    p233 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "00101011001001001100",
            TABLE => "101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p233_in,
            y(0) => p233_out,
            y(1 to 14 - 1) => dummy233
        );


    p234_in <= x(8) & x(17) & x(29) & x(33) & x(70) & x(75) & x(84) & x(90) & x(95) & x(103) & x(117) & x(123) & x(125) & x(126) & x(132) & x(138) & x(242);
    y(234) <= not(p234_out);
    p234 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10011001001100000",
            TABLE => "00101011000000100000001000000000101111110010101100101011000000100010101101000010010000101101010010111101001010110010101101000010011010011001011010010110011010011001011001101001011010011001011001110001000100001111011101110001000100000000000001110001000100000111000100011000111001110111000100011000100011100111000100011000011010011001011010010110011010011001011001101001011010011001011011111110111010001110100010000000011111101110100011101000100000011001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p234_in,
            y(0) => p234_out,
            y(1 to 14 - 1) => dummy234
        );


    p235_in <= x(11) & x(34) & x(52) & x(60) & x(83) & x(89) & x(93) & x(105) & x(112) & x(125) & x(134) & x(135) & x(143) & x(152) & x(188) & x(194) & x(203) & x(204) & x(207) & x(210) & x(216) & x(251);
    y(235) <= not(p235_out);
    p235 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100110110001111000110",
            TABLE => "0001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010011000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010000000000001000000010001000111000001000100011101000111011101111011100010001100000011000100011100001100010001110100011101110011110010110011010010110100110010110011010011001011010010110011010010010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 4,
            B => 6,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p235_in,
            y(0) => p235_out,
            y(1 to 14 - 1) => dummy235
        );


    p236_in <= x(11) & x(27) & x(28) & x(29) & x(40) & x(54) & x(91) & x(93) & x(104) & x(112) & x(118) & x(131) & x(138) & x(179) & x(181) & x(186) & x(240);
    y(236) <= not(p236_out);
    p236 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01000101000101110",
            TABLE => "11010100010000001111110111010100010000000000000011010100010000001101010001000010101111011101010001000010001010111101010001000010100101100110100101101001100101100110100110010110100101100110100111010100010000001111110111010100010000000000000011010100010000001101010001000010101111011101010001000010001010111101010001000010100101100110100101101001100101100110100110010110100101100110100100101011101111110000001000101011001010111011110101000010001010110110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 5,
            B => -8,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p236_in,
            y(0) => p236_out,
            y(1 to 15 - 1) => dummy236
        );


    p237_in <= x(14) & x(24) & x(63) & x(73) & x(77) & x(92) & x(94) & x(114) & x(117) & x(123) & x(136) & x(140) & x(141) & x(154) & x(158) & x(190) & x(227) & x(228) & x(238) & x(253);
    y(237) <= not(p237_out);
    p237 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01100110000100101000",
            TABLE => "010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p237_in,
            y(0) => p237_out,
            y(1 to 14 - 1) => dummy237
        );


    p238_in <= x(5) & x(14) & x(24) & x(37) & x(59) & x(63) & x(73) & x(85) & x(92) & x(175) & x(183) & x(188) & x(189) & x(196) & x(202) & x(240);
    y(238) <= not(p238_out);
    p238 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100101001110010",
            TABLE => "0010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101100001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010011011001000100000101100100010010010010110011010010000000000000000",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p238_in,
            y(0) => p238_out,
            y(1 to 14 - 1) => dummy238
        );


    p239_in <= x(6) & x(7) & x(11) & x(28) & x(51) & x(85) & x(93) & x(100) & x(125) & x(138) & x(140) & x(141) & x(143) & x(163) & x(172) & x(179) & x(182) & x(190) & x(194) & x(199) & x(204) & x(210) & x(225) & x(238) & x(255);
    y(239) <= not(p239_out);
    p239 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1011010100011100111001111",
            TABLE => "0000010001001101000000000000010001001101110111110000010001001101001001000100110110110010001001000100110111011011001001000100110110010110011010010110100110010110011010011001011010010110011010011101010001000000111111011101010001000000000000001101010001000000110101000100001010111101110101000100001000101011110101000100001010010110011010010110100110010110011010011001011010010110011010010001000000000000011100010001000001110001000100001111011101110001000110001000111001110001000110000111000100011000111001110111000110010110011010010110100110010110011010011001011010010110011010010001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010010111",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p239_in,
            y(0) => p239_out,
            y(1 to 14 - 1) => dummy239
        );


    p240_in <= x(15) & x(23) & x(34) & x(58) & x(59) & x(62) & x(83) & x(89) & x(98) & x(113) & x(116) & x(121) & x(125) & x(130) & x(144) & x(147) & x(180) & x(198) & x(202) & x(206) & x(216) & x(219) & x(255);
    y(240) <= not(p240_out);
    p240 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11001100100110011111000",
            TABLE => "00010000000000000111000100010000011100010001000011110111011100010001100010001110011100010001100001110001000110001110011101110001100101100110100101101001100101100110100110010110100101100110100111010100111111010100000011010100010000001101010000000000010000001101010010111101010000101101010001000010110101000010101101000010100101100110100101101001100101100110100110010110100101100110100100010111000000010000000100000000011111110001011100010111000000010001011110000001100000011110100001111110000101110001011110000001100101100110100101101001100101100110100110010110100101100110100110000000111010001110100011111110100000011110100011101000011111101001011001101001011010011001011011111111111111111111111111111111",
            SHIFT => 4,
            B => -5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p240_in,
            y(0) => p240_out,
            y(1 to 14 - 1) => dummy240
        );


    p241_in <= x(0) & x(9) & x(19) & x(25) & x(47) & x(51) & x(55) & x(62) & x(75) & x(76) & x(111) & x(113) & x(133) & x(176) & x(206) & x(228);
    y(241) <= not(p241_out);
    p241 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0111100010000110",
            TABLE => "0000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010011110100011111110100000001110100010000000111010000000000010000000111010000111111010000001111010001000000111101000000101111000000101101001100101101001011001101001100101100110100101101001100101100010101100000010001010110100001001101001100101100000000000000000",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p241_in,
            y(0) => p241_out,
            y(1 to 14 - 1) => dummy241
        );


    p242_in <= x(2) & x(4) & x(10) & x(15) & x(36) & x(61) & x(83) & x(85) & x(89) & x(110) & x(113) & x(144) & x(152) & x(157) & x(162) & x(189) & x(202) & x(212) & x(226) & x(247);
    y(242) <= not(p242_out);
    p242 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10000110101110010100",
            TABLE => "110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 4,
            B => -4,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p242_in,
            y(0) => p242_out,
            y(1 to 14 - 1) => dummy242
        );


    p243_in <= x(23) & x(31) & x(38) & x(56) & x(63) & x(71) & x(81) & x(83) & x(106) & x(160) & x(166) & x(189) & x(196) & x(249);
    y(243) <= not(p243_out);
    p243 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "10100000100000",
            TABLE => "100000001110100000000000100000001110100011111110100000001110100010000001111010000001011110000001111010000111111010000001111010001001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110100010010000",
            SHIFT => 4,
            B => -7,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p243_in,
            y(0) => p243_out,
            y(1 to 13 - 1) => dummy243
        );


    p244_in <= x(5) & x(17) & x(29) & x(32) & x(37) & x(40) & x(48) & x(52) & x(92) & x(95) & x(99) & x(104) & x(112) & x(134) & x(137) & x(138) & x(147) & x(161) & x(164) & x(179) & x(207) & x(232) & x(240) & x(255);
    y(244) <= not(p244_out);
    p244 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100110000000011000011000",
            TABLE => "001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p244_in,
            y(0) => p244_out,
            y(1 to 14 - 1) => dummy244
        );


    p245_in <= x(20) & x(33) & x(36) & x(38) & x(42) & x(49) & x(55) & x(63) & x(72) & x(85) & x(92) & x(111) & x(152) & x(158) & x(164) & x(179) & x(189) & x(193) & x(194) & x(202) & x(206) & x(228) & x(252);
    y(245) <= not(p245_out);
    p245 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "11001001100011011000100",
            TABLE => "00100000000000001011001000100000101100100010000011111011101100100010010001001101101100100010010010110010001001001101101110110010011010011001011010010110011010011001011001101001011010011001011010000000111010001110100011111110000000001000000010000000111010001000000111101000111010000111111000010111100000011000000111101000100101100110100101101001100101100110100110010110100101100110100100000010000000000010101100000010001010110000001010111111001010110100001011010100001010110100001000101011010000101011110100101011100101100110100101101001100101100110100110010110100101100110100111101111100011101000111000001000111001111000111010001110000110000110100110010110100101100110100111111111111111111111111111111111",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p245_in,
            y(0) => p245_out,
            y(1 to 14 - 1) => dummy245
        );


    p246_in <= x(5) & x(11) & x(20) & x(22) & x(29) & x(37) & x(42) & x(46) & x(50) & x(52) & x(56) & x(62) & x(66) & x(69) & x(70) & x(85) & x(94) & x(96) & x(107) & x(111) & x(134) & x(139) & x(142) & x(147) & x(149) & x(154) & x(161) & x(164) & x(179) & x(186) & x(189) & x(248);
    y(246) <= not(p246_out);
    p246 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "01001000011100010101000111110000",
            TABLE => "101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001011111110001011100010111000000010001011100000001000000010000000001111110000101110001011110000001000101111000000110000001111010000110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001110101000100000011111101110101000100000000000000110101000100000011010100010000101011110111010100010000100010101111010100010000101001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001100010010000",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p246_in,
            y(0) => p246_out,
            y(1 to 15 - 1) => dummy246
        );


    p247_in <= x(18) & x(19) & x(25) & x(48) & x(51) & x(66) & x(84) & x(106) & x(117) & x(162) & x(165) & x(166) & x(176) & x(208) & x(209) & x(210) & x(235) & x(239) & x(247);
    y(247) <= not(p247_out);
    p247 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0001110111100110011",
            TABLE => "0111111100010111000101110000000100010111000000010000000100000000011111100001011100010111100000010001011110000001100000011110100001101001100101101001011001101001100101100110100101101001100101100000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010010100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p247_in,
            y(0) => p247_out,
            y(1 to 14 - 1) => dummy247
        );


    p248_in <= x(5) & x(14) & x(27) & x(55) & x(85) & x(92) & x(111) & x(119) & x(157) & x(158) & x(164) & x(168) & x(175) & x(179) & x(181) & x(182) & x(188) & x(193) & x(194) & x(203) & x(206) & x(219) & x(222) & x(246) & x(248);
    y(248) <= not(p248_out);
    p248 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1100000001001100100110101",
            TABLE => "1000000000000000111010001000000011101000100000001111111011101000100000010001011111101000100000011110100010000001011111101110100010010110011010010110100110010110011010011001011010010110011010011110111110001110100011100000100010001110000010000000100000000000111001111000111010001110000110001000111000011000000110000111000101101001100101101001011001101001100101100110100101101001100101100010000000000000101100100010000010110010001000001111101110110010001001000100110110110010001001001011001000100100110110111011001001101001100101101001011001101001100101100110100101101001100101100010000010110010101100101111101100000000001000000010000010110010001001001011001010110010110110110100110100100100001001001011001001101001100101101001011001101001100101100110100101101001100101100111",
            SHIFT => 4,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p248_in,
            y(0) => p248_out,
            y(1 to 14 - 1) => dummy248
        );


    p249_in <= x(6) & x(9) & x(36) & x(40) & x(83) & x(89) & x(94) & x(96) & x(115) & x(141) & x(150) & x(220) & x(234) & x(237) & x(247) & x(249);
    y(249) <= not(p249_out);
    p249 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1110001011101010",
            TABLE => "0000000010000000100000001110100010000000111010001110100011111110000101111000000110000001111010001000000111101000111010000111111001101001100101101001011001101001100101100110100101101001100101100000001000101011000000000000001000101011101111110000001000101011010000100010101111010100010000100010101110111101010000100010101110010110011010010110100110010110011010011001011010010110011010010010000010110010001001001011001001101001100101100000000000000000",
            SHIFT => 5,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p249_in,
            y(0) => p249_out,
            y(1 to 15 - 1) => dummy249
        );


    p250_in <= x(0) & x(3) & x(11) & x(48) & x(55) & x(65) & x(70) & x(117) & x(133) & x(165) & x(168) & x(184) & x(185) & x(186) & x(217) & x(233) & x(235) & x(236);
    y(250) <= not(p250_out);
    p250 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "011000000001100010",
            TABLE => "100000001110100011101000111111100000000010000000100000001110100010000001111010001110100001111110000101111000000110000001111010001001011001101001011010011001011001101001100101101001011001101001111111011101010011010100010000001101010001000000010000000000000010111101110101001101010001000010110101000100001001000010001010110110100110010110100101100110100110010110011010010110100110010110101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => 4,
            B => 3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p250_in,
            y(0) => p250_out,
            y(1 to 14 - 1) => dummy250
        );


    p251_in <= x(7) & x(18) & x(20) & x(30) & x(32) & x(61) & x(63) & x(67) & x(85) & x(87) & x(101) & x(109) & x(113) & x(126) & x(133) & x(148) & x(157) & x(162) & x(174) & x(195) & x(208) & x(212) & x(241) & x(254) & x(255);
    y(251) <= not(p251_out);
    p251 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "1010100000000110111110110",
            TABLE => "0010000010110010000000000010000010110010111110110010000010110010001001001011001001001101001001001011001011011011001001001011001001101001100101101001011001101001100101100110100101101001100101101111111011101000111010001000000011101000100000001000000000000000011111101110100011101000100000011110100010000001100000010001011110010110011010010110100110010110011010011001011010010110011010010001000001110001011100011111011100000000000100000001000001110001000110000111000101110001111001111000111000011000000110000111000110010110011010010110100110010110011010011001011010010110011010010000000000010000000100000111000100010000011100010111000111110111100011100001100000011000011100010001100001110001011100011110011101101001100101101001011001101001100101100110100101101001100101101011",
            SHIFT => 4,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p251_in,
            y(0) => p251_out,
            y(1 to 14 - 1) => dummy251
        );


    p252_in <= x(0) & x(9) & x(19) & x(36) & x(55) & x(63) & x(77) & x(83) & x(85) & x(102) & x(125) & x(126) & x(154) & x(168) & x(171) & x(172) & x(190) & x(193) & x(210) & x(214) & x(224) & x(232) & x(233) & x(238) & x(245) & x(247) & x(254);
    y(252) <= not(p252_out);
    p252 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "100011000110011101011110111",
            TABLE => "011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000101111001011011111111",
            SHIFT => 4,
            B => -2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p252_in,
            y(0) => p252_out,
            y(1 to 14 - 1) => dummy252
        );


    p253_in <= x(3) & x(4) & x(7) & x(10) & x(14) & x(23) & x(24) & x(27) & x(28) & x(31) & x(37) & x(38) & x(51) & x(56) & x(71) & x(73) & x(86) & x(113) & x(121) & x(146) & x(152) & x(179) & x(183) & x(186) & x(188) & x(191) & x(202) & x(205) & x(222) & x(249);
    y(253) <= not(p253_out);
    p253 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "110100111110111000000101010101",
            TABLE => "000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p253_in,
            y(0) => p253_out,
            y(1 to 14 - 1) => dummy253
        );


    p254_in <= x(20) & x(21) & x(33) & x(41) & x(61) & x(66) & x(83) & x(89) & x(102) & x(122) & x(132) & x(137) & x(160) & x(186) & x(197) & x(206) & x(219) & x(225) & x(254);
    y(254) <= not(p254_out);
    p254 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0000101010011001110",
            TABLE => "1111101110110010101100100010000010110010001000000010000000000000110110111011001010110010001001001011001000100100001001000100110101101001100101101001011001101001100101100110100101101001100101100100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100001011100000001000000010000000001111111000101110001011100000001000101111000000110000001111010000111111000010111000101111000000110010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => 2,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p254_in,
            y(0) => p254_out,
            y(1 to 14 - 1) => dummy254
        );


    p255_in <= x(5) & x(16) & x(19) & x(37) & x(61) & x(78) & x(84) & x(102) & x(106) & x(129) & x(141) & x(164) & x(175) & x(181) & x(190) & x(192) & x(205) & x(223) & x(239);
    y(255) <= not(p255_out);
    p255 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "0011001001010001010",
            TABLE => "1000111011101111000010001000111000001000100011100000000000001000100011101110011100011000100011100001100010001110011100010001100010010110011010010110100110010110011010011001011010010110011010010100110100000100000001000000000011011111010011010100110100000100010011010010010000100100101100101101101101001101010011010010010001101001100101101001011001101001100101100110100101101001100101101101111101001101010011010000010001001101000001000000010000000000110110110100110101001101001001000100110100100100001001001011001010010110011010010110100110010110011010011001011010010110011010011011",
            SHIFT => 4,
            B => 5,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p255_in,
            y(0) => p255_out,
            y(1 to 14 - 1) => dummy255
        );



end layer_4;

architecture layer_5 of layer is

    Component perceptron
    Generic (
        WEIGHTS : STD_LOGIC_VECTOR;
        SHIFT : Integer;     -- number of shift (left + or right -)
        B : Integer;          -- bias of batch norm
        BATCH_POSITIVE : Boolean    
    );
    Port ( 
        x : in STD_LOGIC_VECTOR;
        y : out STD_LOGIC_VECTOR
   );
    end component;
    
    -- Signals
    signal p0_in : STD_LOGIC_VECTOR(0 to 81 - 1);
	signal p0_out : STD_LOGIC;
	signal p1_in : STD_LOGIC_VECTOR(0 to 102 - 1);
	signal p1_out : STD_LOGIC;
	signal p2_in : STD_LOGIC_VECTOR(0 to 93 - 1);
	signal p2_out : STD_LOGIC;
	signal p3_in : STD_LOGIC_VECTOR(0 to 87 - 1);
	signal p3_out : STD_LOGIC;
	signal p4_in : STD_LOGIC_VECTOR(0 to 105 - 1);
	signal p4_out : STD_LOGIC;
	signal p5_in : STD_LOGIC_VECTOR(0 to 96 - 1);
	signal p5_out : STD_LOGIC;
	signal p6_in : STD_LOGIC_VECTOR(0 to 92 - 1);
	signal p6_out : STD_LOGIC;
	signal p7_in : STD_LOGIC_VECTOR(0 to 87 - 1);
	signal p7_out : STD_LOGIC;
	signal p8_in : STD_LOGIC_VECTOR(0 to 96 - 1);
	signal p8_out : STD_LOGIC;
	signal p9_in : STD_LOGIC_VECTOR(0 to 112 - 1);
	signal p9_out : STD_LOGIC;
	
    
    -- Dummies
     

begin

    
    p0_in <= x(0) & x(1) & x(4) & x(5) & x(13) & x(20) & x(21) & x(24) & x(28) & x(30) & x(33) & x(37) & x(38) & x(42) & x(47) & x(48) & x(49) & x(51) & x(53) & x(55) & x(58) & x(60) & x(66) & x(70) & x(75) & x(78) & x(80) & x(82) & x(87) & x(88) & x(89) & x(98) & x(100) & x(101) & x(105) & x(112) & x(116) & x(118) & x(119) & x(126) & x(127) & x(128) & x(134) & x(140) & x(141) & x(143) & x(147) & x(148) & x(153) & x(158) & x(161) & x(163) & x(166) & x(176) & x(177) & x(188) & x(191) & x(195) & x(198) & x(199) & x(200) & x(201) & x(205) & x(206) & x(207) & x(213) & x(217) & x(218) & x(225) & x(228) & x(229) & x(231) & x(232) & x(235) & x(241) & x(242) & x(243) & x(245) & x(249) & x(251) & x(254);
    p0 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "",
            TABLE => "000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001010000000000000011010100010000001101010001000000111111011101010001000010001010111101010001000010110101000100001010111101110101000110100110010110100101100110100110010110011010010110100110010110000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110110101000100000001000000000000001111110111010100110101000100000011010100010000100100001000101011101111011101010011010100010000101001011001101001011010011001011001101001100101101001011001101001000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001000101110000000100000001000000000111111100010111000101110000000100010111100000011000000111101000011111100001011100010111100000011001011001101001011010011001011001101001100101101001011001101001000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001110101001001011011111111",
            SHIFT => -3,
            B => -3,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p0_in,
            y => y(0 to 8)
        );


    p1_in <= x(0) & x(3) & x(9) & x(11) & x(19) & x(20) & x(23) & x(25) & x(26) & x(30) & x(32) & x(34) & x(37) & x(39) & x(40) & x(41) & x(42) & x(43) & x(45) & x(46) & x(49) & x(51) & x(54) & x(57) & x(60) & x(63) & x(64) & x(67) & x(68) & x(73) & x(76) & x(77) & x(78) & x(82) & x(83) & x(84) & x(85) & x(89) & x(90) & x(93) & x(94) & x(98) & x(99) & x(100) & x(104) & x(108) & x(109) & x(111) & x(113) & x(114) & x(115) & x(116) & x(117) & x(119) & x(125) & x(126) & x(127) & x(133) & x(136) & x(137) & x(139) & x(141) & x(143) & x(147) & x(148) & x(149) & x(150) & x(151) & x(153) & x(154) & x(155) & x(157) & x(162) & x(170) & x(172) & x(173) & x(174) & x(176) & x(181) & x(182) & x(183) & x(184) & x(194) & x(206) & x(210) & x(212) & x(214) & x(216) & x(218) & x(220) & x(221) & x(229) & x(230) & x(232) & x(233) & x(234) & x(235) & x(238) & x(249) & x(250) & x(252) & x(254);
    p1 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001000101110111111100000001000101110000000100010111000000000000000100010111011111101000000100010111100000010001011111101000100000011001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110000010001000111000000000000010001000111011101111000010001000111000011000100011100111000100011000100011101110011100011000100011100110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111010001000000011111110111010001000000000000000111010001000000011101000100000010111111011101000100000010001011111101000100000010110100110010110100101100110100110010110011010010110100110010110111110111011001010110010001000001011001000100000001000000000000011011011101100101011001000100100101100100010010000100100010011010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => -3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p1_in,
            y => y(9 to 17)
        );


    p2_in <= x(1) & x(6) & x(11) & x(14) & x(15) & x(17) & x(18) & x(20) & x(23) & x(25) & x(26) & x(28) & x(29) & x(31) & x(37) & x(39) & x(42) & x(45) & x(56) & x(58) & x(59) & x(63) & x(64) & x(66) & x(69) & x(72) & x(74) & x(78) & x(85) & x(91) & x(92) & x(93) & x(96) & x(98) & x(101) & x(102) & x(104) & x(111) & x(120) & x(121) & x(122) & x(123) & x(126) & x(127) & x(130) & x(131) & x(135) & x(136) & x(141) & x(142) & x(143) & x(144) & x(148) & x(149) & x(151) & x(153) & x(154) & x(160) & x(164) & x(165) & x(166) & x(169) & x(170) & x(171) & x(173) & x(174) & x(184) & x(186) & x(187) & x(191) & x(192) & x(193) & x(200) & x(201) & x(203) & x(205) & x(207) & x(210) & x(211) & x(214) & x(222) & x(223) & x(225) & x(227) & x(230) & x(232) & x(233) & x(235) & x(245) & x(246) & x(248) & x(251) & x(255);
    p2 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "",
            TABLE => "000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110110101001001011011111111",
            SHIFT => -3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p2_in,
            y => y(18 to 26)
        );


    p3_in <= x(0) & x(2) & x(3) & x(4) & x(5) & x(9) & x(13) & x(15) & x(17) & x(34) & x(36) & x(39) & x(40) & x(41) & x(42) & x(56) & x(58) & x(63) & x(65) & x(66) & x(67) & x(68) & x(69) & x(73) & x(75) & x(78) & x(82) & x(84) & x(85) & x(90) & x(92) & x(97) & x(101) & x(103) & x(106) & x(109) & x(110) & x(112) & x(115) & x(116) & x(117) & x(123) & x(129) & x(137) & x(138) & x(142) & x(149) & x(151) & x(152) & x(157) & x(160) & x(163) & x(167) & x(168) & x(170) & x(176) & x(177) & x(178) & x(182) & x(183) & x(184) & x(186) & x(187) & x(188) & x(189) & x(190) & x(193) & x(195) & x(200) & x(201) & x(203) & x(208) & x(211) & x(217) & x(218) & x(221) & x(223) & x(224) & x(226) & x(231) & x(232) & x(234) & x(237) & x(240) & x(242) & x(251) & x(255);
    p3 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "",
            TABLE => "011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000000010001011100010111011111110000000000000001000000010001011110000001000101110001011101111110111010001000000110000001000101110110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001000000001000000010000000111010001000000011101000111010001111111000010111100000011000000111101000100000011110100011101000011111100110100110010110100101100110100110010110011010010110100110010110001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001011100010110100111111111",
            SHIFT => -3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p3_in,
            y => y(27 to 35)
        );


    p4_in <= x(0) & x(3) & x(4) & x(5) & x(6) & x(7) & x(8) & x(9) & x(11) & x(12) & x(14) & x(15) & x(17) & x(21) & x(23) & x(25) & x(27) & x(28) & x(30) & x(33) & x(35) & x(38) & x(40) & x(43) & x(45) & x(48) & x(57) & x(62) & x(64) & x(66) & x(68) & x(72) & x(73) & x(76) & x(79) & x(80) & x(85) & x(87) & x(89) & x(91) & x(93) & x(95) & x(96) & x(98) & x(111) & x(115) & x(116) & x(117) & x(119) & x(120) & x(121) & x(123) & x(126) & x(127) & x(129) & x(132) & x(136) & x(137) & x(140) & x(142) & x(146) & x(148) & x(150) & x(151) & x(154) & x(155) & x(157) & x(161) & x(162) & x(164) & x(165) & x(175) & x(176) & x(178) & x(181) & x(184) & x(188) & x(191) & x(192) & x(193) & x(194) & x(195) & x(196) & x(197) & x(199) & x(203) & x(205) & x(209) & x(213) & x(217) & x(219) & x(223) & x(224) & x(225) & x(230) & x(232) & x(235) & x(238) & x(240) & x(241) & x(245) & x(246) & x(247) & x(248) & x(252);
    p4 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "",
            TABLE => "101100100010000000100000000000001111101110110010101100100010000010110010001001000010010001001101110110111011001010110010001001001001011001101001011010011001011001101001100101101001011001101001100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001010000001101010000000000010000001101010011111101010000001101010001000010110101000010101101000010110101001011110101000010110101000110100110010110100101100110100110010110011010010110100110010110100000000000000011101000100000001110100010000000111111101110100010000001000101111110100010000001111010001000000101111110111010001001011001101001011010011001011001101001100101101001011001101001000000000000100000001000100011100000100010001110100011101110111101110001000110000001100010001110000110001000111010001110111001111001011001101001011010011001011001101001100101101001011001101001000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110110101001111110101000000110101000100000011010100000000000100000011010100101111010100001011010100010000101101010000101011010000101001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000000100010101100000000000000100010101110111111000000100010101101000010001010111101010001000010001010111011110101000010001010111001011001101001011010011001011001101001100101101001011001101001100011100000100011101111100011100000100000000000100011100000100010001110000110001110011110001110000110000111000110001110000110001001011001101001011010011001011001101001100101101001011001101001000001000100110100000000000001000100110111011111000001000100110100100100010011011011001000100100010011011101101100100100010011011001011001101001011010011001011001101001100101101001011001101001101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001001010110000001000000010000000001011111100101011001010110000001000101011010000100100001011010100101111010010101100101011010000100110100110010110100101100110100110010110011010010110100110010110011100010001000000010000000000001111011101110001011100010001000001110001000110000001100010001110111001110111000101110001000110000110100110010110100101100110100110010110011010010110100110010110001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110000101111001011011111111",
            SHIFT => -3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p4_in,
            y => y(36 to 44)
        );


    p5_in <= x(2) & x(5) & x(6) & x(8) & x(9) & x(11) & x(12) & x(14) & x(15) & x(16) & x(17) & x(21) & x(23) & x(26) & x(28) & x(29) & x(33) & x(36) & x(37) & x(38) & x(39) & x(41) & x(45) & x(47) & x(48) & x(55) & x(58) & x(59) & x(64) & x(65) & x(67) & x(70) & x(71) & x(73) & x(74) & x(75) & x(81) & x(85) & x(87) & x(88) & x(90) & x(93) & x(101) & x(103) & x(106) & x(109) & x(111) & x(112) & x(116) & x(126) & x(128) & x(133) & x(137) & x(138) & x(139) & x(141) & x(143) & x(145) & x(149) & x(150) & x(151) & x(152) & x(153) & x(154) & x(156) & x(162) & x(163) & x(169) & x(170) & x(176) & x(177) & x(181) & x(182) & x(183) & x(190) & x(193) & x(195) & x(201) & x(203) & x(204) & x(206) & x(207) & x(213) & x(215) & x(222) & x(225) & x(226) & x(227) & x(232) & x(234) & x(238) & x(240) & x(242) & x(243) & x(248) & x(253);
    p5 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "",
            TABLE => "001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000100000111000101110001111101110000000000010000000100000111000100011000011100010111000111100111100011100001100000011000011100011001011001101001011010011001011001101001100101101001011001101001101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110000000010001011100000000000000010001011101111111000000010001011110000001000101111110100010000001000101110111111010000001000101110110100110010110100101100110100110010110011010010110100110010110000000100010101100101011101111110000000000000010000000100010101101000010001010110010101110111101110101000100001001000010001010111001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110000101110000000101111111000101110000000100000000000101110000000100010111100000010111111000010111100000011110100000010111100000011001011001101001011010011001011001101001100101101001011001101001001010111011111100000010001010110000001000101011000000000000001000101011101111010100001000101011010000100010101111010100010000100110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001000010001000111010001110111011110000000000001000000010001000111000011000100011101000111011100111011100010001100000011000100011100110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110",
            SHIFT => -3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p5_in,
            y => y(45 to 53)
        );


    p6_in <= x(0) & x(2) & x(3) & x(4) & x(8) & x(11) & x(12) & x(14) & x(15) & x(16) & x(18) & x(19) & x(22) & x(30) & x(37) & x(42) & x(44) & x(45) & x(49) & x(63) & x(67) & x(69) & x(70) & x(73) & x(75) & x(81) & x(84) & x(86) & x(90) & x(95) & x(96) & x(99) & x(101) & x(105) & x(108) & x(109) & x(115) & x(117) & x(121) & x(122) & x(124) & x(130) & x(132) & x(134) & x(140) & x(145) & x(146) & x(147) & x(149) & x(151) & x(155) & x(157) & x(159) & x(164) & x(165) & x(167) & x(168) & x(170) & x(172) & x(173) & x(175) & x(177) & x(178) & x(182) & x(184) & x(187) & x(192) & x(194) & x(198) & x(199) & x(200) & x(209) & x(210) & x(214) & x(216) & x(218) & x(219) & x(220) & x(222) & x(224) & x(227) & x(228) & x(229) & x(230) & x(232) & x(240) & x(244) & x(245) & x(246) & x(249) & x(253) & x(254);
    p6 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "",
            TABLE => "100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110111101110111000101110001000100000111000100010000000100000000000011100111011100010111000100011000011100010001100000011000100011101001011001101001011010011001011001101001100101101001011001101001011100011111011100010000011100010001000001110001000000000001000001110001111001110001100001110001000110000111000110001110000110000110100110010110100101100110100110010110011010010110100110010110100011101110111100001000100011100000100010001110000000000000100010001110111001110001100010001110000110001000111001110001000110001001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001001000000000000010110010001000001011001000100000111110111011001000100100010011011011001000100100101100100010010011011011101100100110100110010110100101100110100110010110011010010110100110010110010011010000010011011111010011010000010000000000010011010000010001001101001001001101101101001101001001001011001001001101001001000110100110010110100101100110100110010110011010010110100110010110101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001001010110000001010111111001010110000001000000000001010110000001000101011010000101011110100101011010000101101010000101011010000100110100110010110100101100110100110010110011010010110100110010110010011011101111100000100010011010000010001001101000000000000010001001101110110110010010001001101001001000100110110110010001001000110100110010110100101100110100110010110011010010110100110010110101100101111101100100000101100100010000010110010000000000010000010110010110110110010010010110010001001001011001001001101001001001001011001101001011010011001011001101001100101101001011001101001101100100010000011111011101100100010000000000000101100100010000010110010001001001101101110110010001001000100110110110010001001001001011001101001011010011001011001101001100101101001011001101001010001100000",
            SHIFT => -3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p6_in,
            y => y(54 to 62)
        );


    p7_in <= x(1) & x(2) & x(3) & x(6) & x(10) & x(14) & x(16) & x(18) & x(19) & x(35) & x(38) & x(40) & x(41) & x(43) & x(46) & x(47) & x(53) & x(54) & x(57) & x(60) & x(65) & x(66) & x(67) & x(69) & x(74) & x(80) & x(81) & x(82) & x(83) & x(86) & x(87) & x(89) & x(91) & x(93) & x(99) & x(103) & x(105) & x(107) & x(115) & x(118) & x(121) & x(123) & x(124) & x(125) & x(127) & x(128) & x(129) & x(131) & x(132) & x(133) & x(134) & x(138) & x(139) & x(143) & x(148) & x(154) & x(159) & x(163) & x(166) & x(172) & x(178) & x(180) & x(185) & x(188) & x(191) & x(194) & x(198) & x(200) & x(202) & x(204) & x(207) & x(216) & x(217) & x(220) & x(223) & x(225) & x(228) & x(231) & x(232) & x(233) & x(237) & x(238) & x(246) & x(247) & x(250) & x(251) & x(252);
    p7 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "",
            TABLE => "001000001011001010110010111110110000000000100000001000001011001000100100101100101011001011011011010011010010010000100100101100100110100110010110100101100110100110010110011010010110100110010110110111110100110101001101000001000100110100000100000001000000000011011011010011010100110100100100010011010010010000100100101100101001011001101001011010011001011001101001100101101001011001101001000001000000000001001101000001000100110100000100110111110100110100100100101100100100110100100100010011010010010011011011010011011001011001101001011010011001011001101001100101101001011001101001001000001011001000000000001000001011001011111011001000001011001000100100101100100100110100100100101100101101101100100100101100100110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001111010001111111010000000111010001000000011101000000000001000000011101000011111101000000111101000100000011110100000010111100000010110100110010110100101100110100110010110011010010110100110010110000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001000100000111000100000000000100000111000111110111000100000111000100011000011100011000111000011000011100011110011100011000011100011001011001101001011010011001011001101001100101101001011001101001000000100000000000101011000000100010101100000010101111110010101101000010110101000010101101000010001010110100001010111101001010111001011001101001011010011001011001101001100101101001011001101001000000000010000000100000101100100010000010110010101100101111101101001101001001000010010010110010001001001011001010110010110110111001011001101001011010011001011001101001100101101001011001101001111111101110100011101000100000001110100010000000100000000000000001111110111010001110100010000001111010001000000110000001000101111001011001101001011010011001011001101001100101101001011001101001000010000000000010001110000010001000111000001000111011111000111000011000011100011000111000011000100011100001100011100111100011100110100110010110100101100110100110010110011010010110100110010110010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110101100101001011011111111",
            SHIFT => -3,
            B => -1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p7_in,
            y => y(63 to 71)
        );


    p8_in <= x(0) & x(1) & x(5) & x(7) & x(8) & x(9) & x(10) & x(11) & x(13) & x(17) & x(18) & x(21) & x(22) & x(28) & x(30) & x(32) & x(36) & x(37) & x(38) & x(39) & x(43) & x(44) & x(46) & x(52) & x(56) & x(57) & x(58) & x(59) & x(60) & x(63) & x(71) & x(73) & x(75) & x(81) & x(84) & x(85) & x(87) & x(88) & x(91) & x(92) & x(95) & x(99) & x(100) & x(101) & x(102) & x(106) & x(111) & x(114) & x(116) & x(120) & x(126) & x(127) & x(129) & x(131) & x(132) & x(135) & x(137) & x(138) & x(141) & x(142) & x(144) & x(146) & x(147) & x(148) & x(151) & x(155) & x(158) & x(160) & x(165) & x(169) & x(170) & x(171) & x(173) & x(177) & x(180) & x(182) & x(183) & x(184) & x(195) & x(196) & x(199) & x(203) & x(207) & x(209) & x(210) & x(211) & x(212) & x(213) & x(220) & x(221) & x(222) & x(226) & x(235) & x(246) & x(249) & x(255);
    p8 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "",
            TABLE => "000000000100000001000000110101000100000011010100110101001111110100101011010000100100001011010100010000101101010011010100101111011001011001101001011010011001011001101001100101101001011001101001010011010000010000000100000000001101111101001101010011010000010001001101001001000010010010110010110110110100110101001101001001000110100110010110100101100110100110010110011010010110100110010110000000000000001000000010001010110000001000101011001010111011111111010100010000100100001000101011010000100010101100101011101111010110100110010110100101100110100110010110011010010110100110010110000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110100011100000100000001000000000001110111110001110100011100000100010001110000110000001100001110001111001111000111010001110000110001001011001101001011010011001011001101001100101101001011001101001000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000000000000010000000100010011010000010001001101010011011101111110110010001001000010010001001101001001000100110101001101110110110110100110010110100101100110100110010110011010010110100110010110000000000000000100000001000101110000000100010111000101110111111111101000100000011000000100010111100000010001011100010111011111101001011001101001011010011001011001101001100101101001011001101001111011111000111010001110000010001000111000001000000010000000000011100111100011101000111000011000100011100001100000011000011100010110100110010110100101100110100110010110011010010110100110010110000000000001000000010000011100010001000001110001011100011111011110001110000110000001100001110001000110000111000101110001111001110110100110010110100101100110100110010110011010010110100110010110101111110010101100101011000000100010101100000010000000100000000010111101001010110010101101000010001010110100001001000010110101001001011001101001011010011001011001101001100101101001011001101001011100010001000011110111011100010001000000000000011100010001000001110001000110001110011101110001000110001000111001110001000110000110100110010110100101100110100110010110011010010110100110010110010000001101010011010100111111010000000001000000010000001101010001000010110101001101010010111101001010110100001001000010110101000110100110010110100101100110100110010110011010010110100110010110000100000000000001110001000100000111000100010000111101110111000100011000100011100111000100011000011100010001100011100111011100011001011001101001011010011001011001101001100101101001011001101001000000010000000000010111000000010001011100000001011111110001011110000001111010000001011110000001000101111000000101111110000101110110100110010110100101100110100110010110011010010110100110010110000001000100110101001101110111110000000000000100000001000100110100100100010011010100110111011011101100100010010000100100010011011001011001101001011010011001011001101001100101101001011001101001",
            SHIFT => -3,
            B => 1,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p8_in,
            y => y(72 to 80)
        );


    p9_in <= x(1) & x(6) & x(9) & x(16) & x(19) & x(21) & x(24) & x(25) & x(30) & x(31) & x(32) & x(33) & x(34) & x(35) & x(36) & x(38) & x(40) & x(42) & x(43) & x(44) & x(47) & x(48) & x(49) & x(52) & x(53) & x(54) & x(56) & x(58) & x(59) & x(60) & x(62) & x(66) & x(68) & x(69) & x(72) & x(74) & x(75) & x(77) & x(78) & x(79) & x(83) & x(84) & x(87) & x(89) & x(91) & x(94) & x(95) & x(96) & x(97) & x(98) & x(100) & x(101) & x(102) & x(105) & x(106) & x(107) & x(108) & x(112) & x(113) & x(117) & x(121) & x(124) & x(125) & x(126) & x(127) & x(128) & x(130) & x(131) & x(132) & x(134) & x(136) & x(137) & x(138) & x(139) & x(153) & x(154) & x(155) & x(161) & x(165) & x(166) & x(167) & x(168) & x(172) & x(173) & x(174) & x(179) & x(182) & x(185) & x(188) & x(190) & x(195) & x(196) & x(199) & x(202) & x(203) & x(205) & x(208) & x(209) & x(213) & x(216) & x(217) & x(218) & x(230) & x(232) & x(233) & x(244) & x(245) & x(246) & x(247) & x(248) & x(250) & x(252);
    p9 : entity work.perceptron(LUT6)
        Generic map (
            WEIGHTS => "",
            TABLE => "1000000011101000111010001111111000000000100000001000000011101000100000011110100011101000011111100001011110000001100000011110100010010110011010010110100110010110011010011001011010010110011010010001011101111111000000010001011100000001000101110000000000000001000101110111111010000001000101111000000100010111111010001000000110010110011010010110100110010110011010011001011010010110011010010100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100001011100000001011111110001011100000001000000000001011100000001000101111000000101111110000101111000000111101000000101111000000110010110011010010110100110010110011010011001011010010110011010010111000100010000111101110111000100010000000000000111000100010000011100010001100011100111011100010001100010001110011100010001100001101001100101101001011001101001100101100110100101101001100101100000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100100110111011111000001000100110100000100010011010000000000000100010011011101101100100100010011010010010001001101101100100010010001101001100101101001011001101001100101100110100101101001100101100100000011010100000000000100000011010100111111010100000011010100010000101101010000101011010000101101010010111101010000101101010001101001100101101001011001101001100101100110100101101001100101100000001000101011001010111011111100000000000000100000001000101011010000100010101100101011101111011101010001000010010000100010101110010110011010010110100110010110011010011001011010010110011010010000000100010111000000000000000100010111011111110000000100010111100000010001011111101000100000010001011101111110100000010001011101101001100101101001011001101001100101100110100101101001100101100000000100010111000101110111111100000000000000010000000100010111100000010001011100010111011111101110100010000001100000010001011101101001100101101001011001101001100101100110100101101001100101100000000000000001000000010001011100000001000101110001011101111111111010001000000110000001000101111000000100010111000101110111111010010110011010010110100110010110011010011001011010010110011010010000010001001101010011011101111100000000000001000000010001001101001001000100110101001101110110111011001000100100001001000100110110010110011010010110100110010110011010011001011010010110011010010100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100000010000000000010011010000010001001101000001001101111101001101001001001011001001001101001001000100110100100100110110110100110110010110011010010110100110010110011010011001011010010110011010010100000011010100110101001111110100000000010000000100000011010100010000101101010011010100101111010010101101000010010000101101010001101001100101101001011001101001100101100110100101101001100101100000000001000000010000001101010001000000110101001101010011111101001010110100001001000010110101000100001011010100110101001011110110010110011010010110100110010110011010011001011010010110011010010100000000000000110101000100000011010100010000001111110111010100010000100010101111010100010000101101010001000010101111011101010001101001100101101001011001101001100101100110100101101001100101100100000011010100010000101101010001101001100101100000000000000000",
            SHIFT => -3,
            B => 0,
            BATCH_POSITIVE => True
        )
        Port map (
            x => p9_in,
            y => y(81 to 89)
        );



end layer_5;
